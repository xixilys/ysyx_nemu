/* verilator lint_off WIDTH */ 
/* verilator lint_off WIDTH */ 
/* verilator lint_off WIDTH */ 
module alu(
  input  [23:0] io_ctrl,
  input  [63:0] io_in1,
  input  [63:0] io_in2,
  output [63:0] io_result,
  output        io_overflow,
  input         io_data_w
);
  wire [5:0] sa = io_in2[5:0]; // @[alu.scala 23:28]
  wire [4:0] sa_for_32bit = io_in2[4:0]; // @[alu.scala 24:30]
  wire [63:0] answer_and = io_in1 & io_in2; // @[alu.scala 26:32]
  wire [63:0] answer_or = io_in1 | io_in2; // @[alu.scala 27:32]
  wire [63:0] answer_xor = io_in1 ^ io_in2; // @[alu.scala 28:32]
  wire [63:0] answer_nor = ~answer_or; // @[alu.scala 29:25]
  wire  answer_slt = $signed(io_in1) < $signed(io_in2); // @[alu.scala 31:43]
  wire  answer_sltu = io_in1 < io_in2; // @[alu.scala 32:36]
  wire [126:0] _GEN_21 = {{63'd0}, io_in1}; // @[alu.scala 33:31]
  wire [126:0] answer_sll = _GEN_21 << sa; // @[alu.scala 33:31]
  wire [63:0] answer_srl = io_in1 >> sa; // @[alu.scala 35:31]
  wire [31:0] answer_srlw = io_in1[31:0] >> sa_for_32bit; // @[alu.scala 36:37]
  wire [63:0] answer_sra = $signed(io_in1) >>> sa; // @[alu.scala 37:46]
  wire [31:0] _answer_sraw_T_1 = io_in1[31:0]; // @[alu.scala 38:38]
  wire [31:0] answer_sraw = $signed(_answer_sraw_T_1) >>> sa_for_32bit; // @[alu.scala 38:62]
  wire [31:0] _answer_lui_T_1 = {io_in2[31:12],12'h0}; // @[Cat.scala 31:58]
  wire [7:0] answer_lui_lo_lo = {_answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],
    _answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31]}; // @[Cat.scala 31:58]
  wire [15:0] answer_lui_lo = {_answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],
    _answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],answer_lui_lo_lo}; // @[Cat.scala 31:58]
  wire [31:0] _answer_lui_T_34 = {_answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],
    _answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],_answer_lui_T_1[31],answer_lui_lo_lo,answer_lui_lo}; // @[Cat.scala 31:58]
  wire [63:0] answer_lui = {_answer_lui_T_34,io_in2[31:12],12'h0}; // @[Cat.scala 31:58]
  wire [64:0] in1_extend = {io_in1[63],io_in1}; // @[Cat.scala 31:58]
  wire [64:0] in2_extend = {io_in2[63],io_in2}; // @[Cat.scala 31:58]
  wire [64:0] answer_add = in1_extend + in2_extend; // @[alu.scala 45:35]
  wire [64:0] answer_sub = in1_extend - in2_extend; // @[alu.scala 46:35]
  wire [23:0] _normal_result_T = {{1'd0}, io_ctrl[23:1]}; // @[alu.scala 49:16]
  wire [23:0] _normal_result_T_3 = {{2'd0}, io_ctrl[23:2]}; // @[alu.scala 50:16]
  wire [23:0] _normal_result_T_6 = {{3'd0}, io_ctrl[23:3]}; // @[alu.scala 51:16]
  wire [23:0] _normal_result_T_9 = {{17'd0}, io_ctrl[23:17]}; // @[alu.scala 52:16]
  wire [23:0] _normal_result_T_12 = {{18'd0}, io_ctrl[23:18]}; // @[alu.scala 53:16]
  wire [23:0] _normal_result_T_15 = {{19'd0}, io_ctrl[23:19]}; // @[alu.scala 54:16]
  wire [23:0] _normal_result_T_18 = {{4'd0}, io_ctrl[23:4]}; // @[alu.scala 55:16]
  wire [23:0] _normal_result_T_20 = {{11'd0}, io_ctrl[23:11]}; // @[alu.scala 56:16]
  wire [23:0] _normal_result_T_22 = {{10'd0}, io_ctrl[23:10]}; // @[alu.scala 57:16]
  wire [23:0] _normal_result_T_24 = {{20'd0}, io_ctrl[23:20]}; // @[alu.scala 58:16]
  wire [23:0] _normal_result_T_26 = {{7'd0}, io_ctrl[23:7]}; // @[alu.scala 59:16]
  wire [23:0] _normal_result_T_28 = {{12'd0}, io_ctrl[23:12]}; // @[alu.scala 60:16]
  wire [23:0] _normal_result_T_30 = {{13'd0}, io_ctrl[23:13]}; // @[alu.scala 61:16]
  wire [23:0] _normal_result_T_32 = {{15'd0}, io_ctrl[23:15]}; // @[alu.scala 62:16]
  wire [63:0] _normal_result_T_34 = io_data_w ? {{32'd0}, answer_sraw} : answer_sra; // @[alu.scala 62:35]
  wire [23:0] _normal_result_T_35 = {{16'd0}, io_ctrl[23:16]}; // @[alu.scala 63:16]
  wire [63:0] _normal_result_T_37 = io_data_w ? {{32'd0}, answer_srlw} : answer_srl; // @[alu.scala 63:35]
  wire [23:0] _normal_result_T_38 = {{14'd0}, io_ctrl[23:14]}; // @[alu.scala 64:16]
  wire [63:0] _normal_result_T_40 = _normal_result_T[0] ? answer_add[63:0] : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_41 = _normal_result_T_3[0] ? answer_add[63:0] : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_42 = _normal_result_T_6[0] ? answer_add[63:0] : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_43 = _normal_result_T_9[0] ? answer_sub[63:0] : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_44 = _normal_result_T_12[0] ? answer_sub[63:0] : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_45 = _normal_result_T_15[0] ? answer_sub[63:0] : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_46 = _normal_result_T_18[0] ? answer_and : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_47 = _normal_result_T_20[0] ? answer_or : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_48 = _normal_result_T_22[0] ? answer_nor : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_49 = _normal_result_T_24[0] ? answer_xor : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_50 = _normal_result_T_26[0] ? answer_lui : 64'h0; // @[Mux.scala 27:73]
  wire [126:0] _normal_result_T_51 = _normal_result_T_28[0] ? answer_sll : 127'h0; // @[Mux.scala 27:73]
  wire  _normal_result_T_52 = _normal_result_T_30[0] & answer_slt; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_53 = _normal_result_T_32[0] ? _normal_result_T_34 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_54 = _normal_result_T_35[0] ? _normal_result_T_37 : 64'h0; // @[Mux.scala 27:73]
  wire  _normal_result_T_55 = _normal_result_T_38[0] & answer_sltu; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_56 = _normal_result_T_40 | _normal_result_T_41; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_57 = _normal_result_T_56 | _normal_result_T_42; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_58 = _normal_result_T_57 | _normal_result_T_43; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_59 = _normal_result_T_58 | _normal_result_T_44; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_60 = _normal_result_T_59 | _normal_result_T_45; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_61 = _normal_result_T_60 | _normal_result_T_46; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_62 = _normal_result_T_61 | _normal_result_T_47; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_63 = _normal_result_T_62 | _normal_result_T_48; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_64 = _normal_result_T_63 | _normal_result_T_49; // @[Mux.scala 27:73]
  wire [63:0] _normal_result_T_65 = _normal_result_T_64 | _normal_result_T_50; // @[Mux.scala 27:73]
  wire [126:0] _GEN_16 = {{63'd0}, _normal_result_T_65}; // @[Mux.scala 27:73]
  wire [126:0] _normal_result_T_66 = _GEN_16 | _normal_result_T_51; // @[Mux.scala 27:73]
  wire [126:0] _GEN_17 = {{126'd0}, _normal_result_T_52}; // @[Mux.scala 27:73]
  wire [126:0] _normal_result_T_67 = _normal_result_T_66 | _GEN_17; // @[Mux.scala 27:73]
  wire [126:0] _GEN_18 = {{63'd0}, _normal_result_T_53}; // @[Mux.scala 27:73]
  wire [126:0] _normal_result_T_68 = _normal_result_T_67 | _GEN_18; // @[Mux.scala 27:73]
  wire [126:0] _GEN_19 = {{63'd0}, _normal_result_T_54}; // @[Mux.scala 27:73]
  wire [126:0] _normal_result_T_69 = _normal_result_T_68 | _GEN_19; // @[Mux.scala 27:73]
  wire [126:0] _GEN_20 = {{126'd0}, _normal_result_T_55}; // @[Mux.scala 27:73]
  wire [126:0] normal_result = _normal_result_T_69 | _GEN_20; // @[Mux.scala 27:73]
  wire [7:0] io_result_lo_lo = {normal_result[31],normal_result[31],normal_result[31],normal_result[31],normal_result[31
    ],normal_result[31],normal_result[31],normal_result[31]}; // @[Cat.scala 31:58]
  wire [15:0] io_result_lo = {normal_result[31],normal_result[31],normal_result[31],normal_result[31],normal_result[31],
    normal_result[31],normal_result[31],normal_result[31],io_result_lo_lo}; // @[Cat.scala 31:58]
  wire [31:0] _io_result_T_33 = {normal_result[31],normal_result[31],normal_result[31],normal_result[31],normal_result[
    31],normal_result[31],normal_result[31],normal_result[31],io_result_lo_lo,io_result_lo}; // @[Cat.scala 31:58]
  wire [63:0] _io_result_T_35 = {_io_result_T_33,normal_result[31:0]}; // @[Cat.scala 31:58]
  wire [126:0] _io_result_T_36 = io_data_w ? {{63'd0}, _io_result_T_35} : normal_result; // @[alu.scala 66:21]
  assign io_result = _io_result_T_36[63:0]; // @[alu.scala 66:15]
  assign io_overflow = _normal_result_T_3[0] & answer_add[64] != answer_add[63] | _normal_result_T_12[0] & answer_sub[64
    ] != answer_sub[63]; // @[alu.scala 67:101]
endmodule
module br(
  input         reset,
  input  [63:0] io_r1,
  input  [63:0] io_r2,
  input  [5:0]  io_branch,
  output        io_exe
);
  wire  _result_T = io_r1 >= io_r2; // @[br.scala 24:38]
  wire  _result_T_1 = io_r1 < io_r2; // @[br.scala 25:37]
  wire  _result_T_4 = $signed(io_r1) >= $signed(io_r2); // @[br.scala 26:37]
  wire  _result_T_7 = $signed(io_r1) < $signed(io_r2); // @[br.scala 27:37]
  wire  _result_T_8 = io_r1 != io_r2; // @[br.scala 28:30]
  wire  _result_T_9 = io_r1 == io_r2; // @[br.scala 29:30]
  wire [5:0] result = {_result_T,_result_T_1,_result_T_4,_result_T_7,_result_T_8,_result_T_9}; // @[Cat.scala 31:58]
  wire [5:0] _io_exe_T_4 = result & io_branch; // @[br.scala 30:57]
  assign io_exe = ~reset & _io_exe_T_4 != 6'h0; // @[br.scala 30:45]
endmodule
module cfu(
  input         reset,
  input         io_Inst_Fifo_Empty,
  input         io_dmem_calD,
  input         io_BranchD_Flag,
  input         io_JRD,
  input         io_CanBranchD,
  input         io_DivPendingE,
  input         io_DataPendingM,
  input         io_InException,
  input  [4:0]  io_WriteRegE,
  input         io_RegWriteE,
  input         io_csrToRegE,
  input  [4:0]  io_WriteRegM,
  input         io_MemToRegM,
  input         io_RegWriteM,
  input         io_csrWriteM,
  input  [4:0]  io_WriteRegM2,
  input         io_MemToRegM2,
  input         io_RegWriteM2,
  input         io_csrWriteM2,
  input  [4:0]  io_WriteRegW,
  input         io_RegWriteW,
  input  [11:0] io_ReadcsrAddrE,
  input  [11:0] io_WritecsrAddrM,
  input  [11:0] io_WritecsrAddrM2,
  input  [4:0]  io_R2D,
  input  [4:0]  io_R1D,
  input  [4:0]  io_R2E,
  input  [4:0]  io_R1E,
  output        io_StallF,
  output        io_StallD,
  output        io_StallE,
  output        io_StallM,
  output        io_StallM2,
  output        io_StallW,
  output        io_FlushD,
  output        io_FlushE,
  output        io_FlushM,
  output        io_FlushM2,
  output        io_FlushW,
  output [1:0]  io_Forward1E,
  output [1:0]  io_Forward2E,
  output [1:0]  io_Forward1D,
  output [1:0]  io_Forward2D,
  output [1:0]  io_ForwardcsrE
);
  wire  _io_Forward2D_T_3 = io_R2D == io_WriteRegM & io_RegWriteM; // @[cfu.scala 94:73]
  wire  _io_Forward2D_T_5 = ~io_MemToRegM; // @[cfu.scala 94:99]
  wire  _io_Forward2D_T_9 = io_R2D == io_WriteRegM2 & io_RegWriteM2; // @[cfu.scala 95:34]
  wire  _io_Forward2D_T_11 = ~io_MemToRegM2; // @[cfu.scala 95:61]
  wire  _io_Forward2D_T_12 = io_R2D == io_WriteRegM2 & io_RegWriteM2 & ~io_MemToRegM2; // @[cfu.scala 95:58]
  wire [1:0] _io_Forward2D_T_13 = _io_Forward2D_T_12 ? 2'h2 : 2'h0; // @[cfu.scala 94:131]
  wire [1:0] _io_Forward2D_T_14 = io_R2D == io_WriteRegM & io_RegWriteM & ~io_MemToRegM ? 2'h1 : _io_Forward2D_T_13; // @[cfu.scala 94:48]
  wire  _io_Forward1D_T_3 = io_R1D == io_WriteRegM & io_RegWriteM; // @[cfu.scala 96:73]
  wire  _io_Forward1D_T_9 = io_R1D == io_WriteRegM2 & io_RegWriteM2; // @[cfu.scala 97:34]
  wire  _io_Forward1D_T_12 = io_R1D == io_WriteRegM2 & io_RegWriteM2 & _io_Forward2D_T_11; // @[cfu.scala 97:58]
  wire [1:0] _io_Forward1D_T_13 = _io_Forward1D_T_12 ? 2'h2 : 2'h0; // @[cfu.scala 96:131]
  wire [1:0] _io_Forward1D_T_14 = io_R1D == io_WriteRegM & io_RegWriteM & _io_Forward2D_T_5 ? 2'h1 : _io_Forward1D_T_13; // @[cfu.scala 96:48]
  wire  _io_Forward2E_T_3 = io_R2E == io_WriteRegM & io_RegWriteM; // @[cfu.scala 103:34]
  wire  _io_Forward2E_T_6 = io_R2E == io_WriteRegM & io_RegWriteM & _io_Forward2D_T_5; // @[cfu.scala 103:57]
  wire  _io_Forward2E_T_9 = io_R2E == io_WriteRegM2 & io_RegWriteM2; // @[cfu.scala 104:35]
  wire  _io_Forward2E_T_12 = io_R2E == io_WriteRegM2 & io_RegWriteM2 & _io_Forward2D_T_11; // @[cfu.scala 104:59]
  wire  _io_Forward2E_T_15 = io_R2E == io_WriteRegW & io_RegWriteW; // @[cfu.scala 105:34]
  wire [1:0] _io_Forward2E_T_17 = _io_Forward2E_T_12 ? 2'h3 : {{1'd0}, _io_Forward2E_T_15}; // @[Mux.scala 101:16]
  wire [1:0] _io_Forward2E_T_18 = _io_Forward2E_T_6 ? 2'h2 : _io_Forward2E_T_17; // @[Mux.scala 101:16]
  wire  _io_Forward1E_T_3 = io_R1E == io_WriteRegM & io_RegWriteM; // @[cfu.scala 110:34]
  wire  _io_Forward1E_T_6 = io_R1E == io_WriteRegM & io_RegWriteM & _io_Forward2D_T_5; // @[cfu.scala 110:57]
  wire  _io_Forward1E_T_9 = io_R1E == io_WriteRegM2 & io_RegWriteM2; // @[cfu.scala 111:35]
  wire  _io_Forward1E_T_12 = io_R1E == io_WriteRegM2 & io_RegWriteM2 & _io_Forward2D_T_11; // @[cfu.scala 111:59]
  wire  _io_Forward1E_T_15 = io_R1E == io_WriteRegW & io_RegWriteW; // @[cfu.scala 112:34]
  wire [1:0] _io_Forward1E_T_17 = _io_Forward1E_T_12 ? 2'h3 : {{1'd0}, _io_Forward1E_T_15}; // @[Mux.scala 101:16]
  wire [1:0] _io_Forward1E_T_18 = _io_Forward1E_T_6 ? 2'h2 : _io_Forward1E_T_17; // @[Mux.scala 101:16]
  wire  _io_ForwardcsrE_T_3 = io_ReadcsrAddrE == io_WritecsrAddrM & io_csrWriteM; // @[cfu.scala 118:59]
  wire  _io_ForwardcsrE_T_6 = io_ReadcsrAddrE == io_WritecsrAddrM2 & io_csrWriteM2; // @[cfu.scala 119:60]
  wire [1:0] _io_ForwardcsrE_T_7 = _io_ForwardcsrE_T_6 ? 2'h2 : 2'h0; // @[Mux.scala 101:16]
  wire [1:0] _io_ForwardcsrE_T_8 = _io_ForwardcsrE_T_3 ? 2'h1 : _io_ForwardcsrE_T_7; // @[Mux.scala 101:16]
  wire  _br_Stall_T_5 = io_WriteRegE == io_R1D; // @[cfu.scala 125:75]
  wire  _br_Stall_T_10 = io_WriteRegM == io_R1D; // @[cfu.scala 126:74]
  wire  _br_Stall_T_12 = io_MemToRegM & (io_WriteRegM == io_R2D | io_WriteRegM == io_R1D); // @[cfu.scala 126:30]
  wire  _br_Stall_T_13 = io_RegWriteE & (io_WriteRegE == io_R2D | io_WriteRegE == io_R1D) | _br_Stall_T_12; // @[cfu.scala 125:88]
  wire  _br_Stall_T_16 = io_WriteRegM2 == io_R1D; // @[cfu.scala 127:77]
  wire  _br_Stall_T_18 = io_MemToRegM2 & (io_WriteRegM2 == io_R2D | io_WriteRegM2 == io_R1D); // @[cfu.scala 127:31]
  wire  _br_Stall_T_19 = _br_Stall_T_13 | _br_Stall_T_18; // @[cfu.scala 126:87]
  wire  _br_Stall_T_20 = io_CanBranchD & io_BranchD_Flag & _br_Stall_T_19; // @[cfu.scala 124:71]
  wire  _br_Stall_T_22 = ~io_InException; // @[cfu.scala 127:95]
  wire  br_Stall = _br_Stall_T_20 & ~io_InException; // @[cfu.scala 127:92]
  wire  _jr_Stall_T_8 = io_MemToRegM & _br_Stall_T_10; // @[cfu.scala 130:30]
  wire  _jr_Stall_T_9 = io_RegWriteE & _br_Stall_T_5 | _jr_Stall_T_8; // @[cfu.scala 129:61]
  wire  _jr_Stall_T_12 = io_MemToRegM2 & _br_Stall_T_16; // @[cfu.scala 131:31]
  wire  _jr_Stall_T_13 = _jr_Stall_T_9 | _jr_Stall_T_12; // @[cfu.scala 130:62]
  wire  _jr_Stall_T_14 = (io_JRD | io_dmem_calD) & _jr_Stall_T_13; // @[cfu.scala 128:60]
  wire  dmem_addr_cal_Stall = _jr_Stall_T_14 & _br_Stall_T_22; // @[cfu.scala 131:65]
  wire  _mem2regM_Stall_T_9 = _io_Forward1E_T_3 & io_MemToRegM; // @[cfu.scala 142:87]
  wire  _mem2regM_Stall_T_10 = _io_Forward2E_T_3 & io_MemToRegM | _mem2regM_Stall_T_9; // @[cfu.scala 141:120]
  wire  _mem2regM_Stall_T_15 = _io_Forward2D_T_3 & io_MemToRegM; // @[cfu.scala 143:87]
  wire  _mem2regM_Stall_T_16 = _mem2regM_Stall_T_10 | _mem2regM_Stall_T_15; // @[cfu.scala 142:111]
  wire  _mem2regM_Stall_T_21 = _io_Forward1D_T_3 & io_MemToRegM; // @[cfu.scala 144:87]
  wire  _mem2regM_Stall_T_22 = _mem2regM_Stall_T_16 | _mem2regM_Stall_T_21; // @[cfu.scala 143:111]
  wire  _mem2regM_Stall_T_27 = _io_Forward2E_T_9 & io_MemToRegM2; // @[cfu.scala 145:89]
  wire  _mem2regM_Stall_T_28 = _mem2regM_Stall_T_22 | _mem2regM_Stall_T_27; // @[cfu.scala 144:111]
  wire  _mem2regM_Stall_T_33 = _io_Forward1E_T_9 & io_MemToRegM2; // @[cfu.scala 146:89]
  wire  _mem2regM_Stall_T_34 = _mem2regM_Stall_T_28 | _mem2regM_Stall_T_33; // @[cfu.scala 145:114]
  wire  _mem2regM_Stall_T_39 = _io_Forward2D_T_9 & io_MemToRegM2; // @[cfu.scala 147:89]
  wire  _mem2regM_Stall_T_40 = _mem2regM_Stall_T_34 | _mem2regM_Stall_T_39; // @[cfu.scala 146:114]
  wire  _mem2regM_Stall_T_45 = _io_Forward1D_T_9 & io_MemToRegM2; // @[cfu.scala 148:89]
  wire  mem2regM_Stall = _mem2regM_Stall_T_40 | _mem2regM_Stall_T_45; // @[cfu.scala 147:114]
  wire  _has_Stall_T = br_Stall | dmem_addr_cal_Stall; // @[cfu.scala 155:44]
  wire  _io_StallF_T_5 = _has_Stall_T | io_DivPendingE | io_DataPendingM | mem2regM_Stall; // @[cfu.scala 160:133]
  wire  _io_StallM_T_1 = ~io_DataPendingM; // @[cfu.scala 163:39]
  assign io_StallF = reset | ~(_has_Stall_T | io_DivPendingE | io_DataPendingM | mem2regM_Stall | io_Inst_Fifo_Empty); // @[cfu.scala 160:21]
  assign io_StallD = reset | ~_io_StallF_T_5; // @[cfu.scala 161:21]
  assign io_StallE = reset | ~(io_DivPendingE | io_DataPendingM | mem2regM_Stall); // @[cfu.scala 162:21]
  assign io_StallM = reset | ~io_DataPendingM; // @[cfu.scala 163:21]
  assign io_StallM2 = reset | _io_StallM_T_1; // @[cfu.scala 164:22]
  assign io_StallW = reset | _io_StallM_T_1; // @[cfu.scala 165:21]
  assign io_FlushD = reset ? 1'h0 : io_InException; // @[cfu.scala 167:21]
  assign io_FlushE = reset ? 1'h0 : io_StallE & _has_Stall_T | io_InException; // @[cfu.scala 168:21]
  assign io_FlushM = reset ? 1'h0 : io_StallM & (io_DivPendingE | mem2regM_Stall) | io_InException; // @[cfu.scala 169:21]
  assign io_FlushM2 = reset ? 1'h0 : io_InException; // @[cfu.scala 170:22]
  assign io_FlushW = reset ? 1'h0 : io_StallW & (io_DataPendingM | io_InException); // @[cfu.scala 171:21]
  assign io_Forward1E = io_R1E == 5'h0 ? 2'h0 : _io_Forward1E_T_18; // @[cfu.scala 109:24]
  assign io_Forward2E = io_R2E == 5'h0 ? 2'h0 : _io_Forward2E_T_18; // @[cfu.scala 102:24]
  assign io_Forward1D = io_R1D == 5'h0 ? 2'h0 : _io_Forward1D_T_14; // @[cfu.scala 96:24]
  assign io_Forward2D = io_R2D == 5'h0 ? 2'h0 : _io_Forward2D_T_14; // @[cfu.scala 94:24]
  assign io_ForwardcsrE = io_csrToRegE ? _io_ForwardcsrE_T_8 : 2'h0; // @[cfu.scala 117:26]
endmodule
module csr(
  input         clock,
  input         reset,
  input  [11:0] io_csr_read_addr,
  input  [11:0] io_csr_write_addr,
  input  [63:0] io_csr_write_data,
  input         io_csr_write_en,
  input  [63:0] io_pc,
  input  [31:0] io_exception_type_i,
  output [63:0] io_return_pc,
  output        io_exception,
  output [63:0] io_csr_read_data,
  output        io_icache_tags_flush,
  input         io_int_type_timer,
  output        io_Int_able,
  output        io_int_type_able_timer
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] csr_cause; // @[csr.scala 59:28]
  reg [63:0] csr_status; // @[csr.scala 60:25]
  wire  _csr_status_to_be_T_3 = io_csr_write_en & io_csr_write_addr == 12'h300; // @[csr.scala 175:33]
  wire  csr_status_to_vec_63 = csr_status[63]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_62 = csr_status[62]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_61 = csr_status[61]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_60 = csr_status[60]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_59 = csr_status[59]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_58 = csr_status[58]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_57 = csr_status[57]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_56 = csr_status[56]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_55 = csr_status[55]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_54 = csr_status[54]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_53 = csr_status[53]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_52 = csr_status[52]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_51 = csr_status[51]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_50 = csr_status[50]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_49 = csr_status[49]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_48 = csr_status[48]; // @[csr.scala 167:28]
  wire [7:0] csr_status_to_be_hi_hi_lo = {csr_status_to_vec_55,csr_status_to_vec_54,csr_status_to_vec_53,
    csr_status_to_vec_52,csr_status_to_vec_51,csr_status_to_vec_50,csr_status_to_vec_49,csr_status_to_vec_48}; // @[csr.scala 174:53]
  wire  csr_status_to_vec_47 = csr_status[47]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_46 = csr_status[46]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_45 = csr_status[45]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_44 = csr_status[44]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_43 = csr_status[43]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_42 = csr_status[42]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_41 = csr_status[41]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_40 = csr_status[40]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_39 = csr_status[39]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_38 = csr_status[38]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_37 = csr_status[37]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_36 = csr_status[36]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_35 = csr_status[35]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_34 = csr_status[34]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_33 = csr_status[33]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_32 = csr_status[32]; // @[csr.scala 167:28]
  wire [7:0] csr_status_to_be_hi_lo_lo = {csr_status_to_vec_39,csr_status_to_vec_38,csr_status_to_vec_37,
    csr_status_to_vec_36,csr_status_to_vec_35,csr_status_to_vec_34,csr_status_to_vec_33,csr_status_to_vec_32}; // @[csr.scala 174:53]
  wire [15:0] csr_status_to_be_hi_lo = {csr_status_to_vec_47,csr_status_to_vec_46,csr_status_to_vec_45,
    csr_status_to_vec_44,csr_status_to_vec_43,csr_status_to_vec_42,csr_status_to_vec_41,csr_status_to_vec_40,
    csr_status_to_be_hi_lo_lo}; // @[csr.scala 174:53]
  wire [31:0] csr_status_to_be_hi = {csr_status_to_vec_63,csr_status_to_vec_62,csr_status_to_vec_61,csr_status_to_vec_60
    ,csr_status_to_vec_59,csr_status_to_vec_58,csr_status_to_vec_57,csr_status_to_vec_56,csr_status_to_be_hi_hi_lo,
    csr_status_to_be_hi_lo}; // @[csr.scala 174:53]
  wire  csr_status_to_vec_31 = csr_status[31]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_30 = csr_status[30]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_29 = csr_status[29]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_28 = csr_status[28]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_27 = csr_status[27]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_26 = csr_status[26]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_25 = csr_status[25]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_24 = csr_status[24]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_23 = csr_status[23]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_22 = csr_status[22]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_21 = csr_status[21]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_20 = csr_status[20]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_19 = csr_status[19]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_18 = csr_status[18]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_17 = csr_status[17]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_16 = csr_status[16]; // @[csr.scala 167:28]
  wire [7:0] csr_status_to_be_lo_hi_lo = {csr_status_to_vec_23,csr_status_to_vec_22,csr_status_to_vec_21,
    csr_status_to_vec_20,csr_status_to_vec_19,csr_status_to_vec_18,csr_status_to_vec_17,csr_status_to_vec_16}; // @[csr.scala 174:53]
  wire  csr_status_to_vec_15 = csr_status[15]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_14 = csr_status[14]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_13 = csr_status[13]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_12 = csr_status[12]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_11 = csr_status[11]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_10 = csr_status[10]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_9 = csr_status[9]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_8 = csr_status[8]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_7 = csr_status[7]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_6 = csr_status[6]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_5 = csr_status[5]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_4 = csr_status[4]; // @[csr.scala 167:28]
  reg [63:0] csr_mie; // @[csr.scala 71:28]
  wire  csr_status_to_vec_3 = csr_status[3]; // @[csr.scala 165:54]
  wire  csr_status_to_vec_2 = csr_status[2]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_1 = csr_status[1]; // @[csr.scala 167:28]
  wire  csr_status_to_vec_0 = csr_status[0]; // @[csr.scala 167:28]
  wire [7:0] csr_status_to_be_lo_lo_lo = {csr_status_to_vec_7,csr_status_to_vec_6,csr_status_to_vec_5,
    csr_status_to_vec_4,csr_status_to_vec_3,csr_status_to_vec_2,csr_status_to_vec_1,csr_status_to_vec_0}; // @[csr.scala 174:53]
  wire [15:0] csr_status_to_be_lo_lo = {csr_status_to_vec_15,csr_status_to_vec_14,csr_status_to_vec_13,
    csr_status_to_vec_12,csr_status_to_vec_11,csr_status_to_vec_10,csr_status_to_vec_9,csr_status_to_vec_8,
    csr_status_to_be_lo_lo_lo}; // @[csr.scala 174:53]
  wire [31:0] csr_status_to_be_lo = {csr_status_to_vec_31,csr_status_to_vec_30,csr_status_to_vec_29,csr_status_to_vec_28
    ,csr_status_to_vec_27,csr_status_to_vec_26,csr_status_to_vec_25,csr_status_to_vec_24,csr_status_to_be_lo_hi_lo,
    csr_status_to_be_lo_lo}; // @[csr.scala 174:53]
  wire [63:0] _csr_status_to_be_T = {csr_status_to_be_hi,csr_status_to_be_lo}; // @[csr.scala 174:53]
  reg [63:0] csr_epc; // @[csr.scala 63:26]
  reg [63:0] csr_mtvec; // @[csr.scala 64:28]
  reg [63:0] csr_mip; // @[csr.scala 72:28]
  wire [31:0] exception_type = {io_exception_type_i[31:1],1'h0}; // @[Cat.scala 31:58]
  wire [31:0] _commit_exception_T_2 = {{24'd0}, exception_type[31:24]}; // @[csr.scala 90:76]
  wire  commit_exception = exception_type[30:0] != 31'h0 & ~_commit_exception_T_2[0]; // @[csr.scala 90:58]
  wire [31:0] _commit_eret_T_1 = {{20'd0}, exception_type[31:20]}; // @[csr.scala 91:65]
  wire  commit_eret = exception_type[31] & ~_commit_eret_T_1[0]; // @[csr.scala 91:47]
  wire [63:0] _csr_read_data_Wire_T_1 = 12'h341 == io_csr_read_addr ? csr_epc : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _csr_read_data_Wire_T_3 = 12'h342 == io_csr_read_addr ? csr_cause : _csr_read_data_Wire_T_1; // @[Mux.scala 81:58]
  wire [63:0] _csr_read_data_Wire_T_5 = 12'h305 == io_csr_read_addr ? csr_mtvec : _csr_read_data_Wire_T_3; // @[Mux.scala 81:58]
  wire [63:0] _csr_read_data_Wire_T_7 = 12'h300 == io_csr_read_addr ? csr_status : _csr_read_data_Wire_T_5; // @[Mux.scala 81:58]
  wire [63:0] _csr_read_data_Wire_T_9 = 12'h344 == io_csr_read_addr ? csr_mip : _csr_read_data_Wire_T_7; // @[Mux.scala 81:58]
  wire [63:0] csr_read_data_Wire = 12'h304 == io_csr_read_addr ? csr_mie : _csr_read_data_Wire_T_9; // @[Mux.scala 81:58]
  wire [63:0] _io_return_pc_T_2 = io_pc + 64'h4; // @[csr.scala 106:38]
  wire [63:0] _io_return_pc_T_3 = _commit_exception_T_2[0] ? _io_return_pc_T_2 : csr_mtvec; // @[Mux.scala 101:16]
  wire [31:0] _cause_exccode_T_3 = {{8'd0}, exception_type[31:8]}; // @[csr.scala 119:23]
  wire [63:0] _cause_exccode_T_5 = exception_type[0] ? 64'h8000000000000011 : 64'h0; // @[Mux.scala 27:73]
  wire [3:0] _cause_exccode_T_6 = _cause_exccode_T_3[0] ? 4'hb : 4'h0; // @[Mux.scala 27:73]
  wire [63:0] _GEN_4 = {{60'd0}, _cause_exccode_T_6}; // @[Mux.scala 27:73]
  wire [63:0] cause_exccode = _cause_exccode_T_5 | _GEN_4; // @[Mux.scala 27:73]
  wire  _csr_epc_T_3 = io_csr_write_en & io_csr_write_addr == 12'h341; // @[csr.scala 172:32]
  wire  _csr_mtvec_T_2 = io_csr_write_en & io_csr_write_addr == 12'h305; // @[csr.scala 178:33]
  wire  _csr_cause_T_2 = io_csr_write_en & io_csr_write_addr == 12'h342; // @[csr.scala 181:33]
  wire  _csr_mie_T_2 = io_csr_write_en & io_csr_write_addr == 12'h304; // @[csr.scala 186:33]
  wire [63:0] _csr_mip_T = {32'h0,16'h0,8'h0,io_int_type_timer,1'h0,2'h0,4'h0}; // @[csr.scala 195:42]
  wire  _csr_mip_T_3 = io_csr_write_en & io_csr_write_addr == 12'h344; // @[csr.scala 196:33]
  assign io_return_pc = commit_eret ? csr_epc : _io_return_pc_T_3; // @[Mux.scala 101:16]
  assign io_exception = commit_exception | commit_eret; // @[csr.scala 93:43]
  assign io_csr_read_data = reset ? 64'h0 : csr_read_data_Wire; // @[csr.scala 100:29]
  assign io_icache_tags_flush = _commit_exception_T_2[0]; // @[csr.scala 92:40]
  assign io_Int_able = csr_status[3]; // @[csr.scala 159:30]
  assign io_int_type_able_timer = csr_mie[7]; // @[csr.scala 189:38]
  always @(posedge clock) begin
    if (reset) begin // @[csr.scala 62:22]
      csr_status <= 64'ha00001800;
    end else if (_csr_status_to_be_T_3) begin // @[Mux.scala 101:16]
      csr_status <= io_csr_write_data;
    end else begin
      csr_status <= _csr_status_to_be_T;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Mux.scala 101:16]
      csr_cause <= 64'h400000;
    end else if (_csr_cause_T_2) begin // @[Mux.scala 101:16]
      csr_cause <= io_csr_write_data;
    end else if (commit_exception) begin
      csr_cause <= cause_exccode;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Mux.scala 101:16]
      csr_mie <= 64'h0;
    end else if (_csr_mie_T_2) begin
      csr_mie <= io_csr_write_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Mux.scala 101:16]
      csr_epc <= 64'h0;
    end else if (commit_exception) begin // @[Mux.scala 101:16]
      csr_epc <= io_pc;
    end else if (_csr_epc_T_3) begin
      csr_epc <= io_csr_write_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Mux.scala 101:16]
      csr_mtvec <= 64'h0;
    end else if (_csr_mtvec_T_2) begin
      csr_mtvec <= io_csr_write_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Mux.scala 101:16]
      csr_mip <= 64'h0;
    end else if (_csr_mip_T_3) begin
      csr_mip <= io_csr_write_data;
    end else begin
      csr_mip <= _csr_mip_T;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  csr_cause = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  csr_status = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  csr_mie = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  csr_epc = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  csr_mtvec = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  csr_mip = _RAND_5[63:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    csr_cause = 64'h400000;
  end
  if (reset) begin
    csr_mie = 64'h0;
  end
  if (reset) begin
    csr_epc = 64'h0;
  end
  if (reset) begin
    csr_mtvec = 64'h0;
  end
  if (reset) begin
    csr_mip = 64'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module cu(
  input  [31:0] io1_InstrD,
  output        io1_BadInstrD,
  output        io1_SysCallD,
  output        io1_EretD,
  output        io1_dmem_addr_cal,
  output        io_RegWriteD,
  output        io_MemToRegD,
  output        io_MemWriteD,
  output [23:0] io_ALUCtrlD,
  output [1:0]  io_ALUSrcD_0,
  output [1:0]  io_ALUSrcD_1,
  output [4:0]  io_RegDstD,
  output        io_LinkD,
  output        io_csrWriteD,
  output        io_csrToRegD,
  output        io_LoadUnsignedD,
  output [1:0]  io_MemWidthD,
  output [63:0] io_ImmD,
  output        io_ebreakD,
  output        io_data_wD,
  output [23:0] io_muldiv_control,
  output        io_muldiv_cal,
  output        io_alu_cal,
  output [5:0]  io_csr_control,
  output        io_csr_Imm,
  output        io_fence_i_control
);
  wire [6:0] OpD = io1_InstrD[6:0]; // @[cu.scala 63:25]
  wire [2:0] Funct3D = io1_InstrD[14:12]; // @[cu.scala 64:29]
  wire [6:0] Funct7D = io1_InstrD[31:25]; // @[cu.scala 65:29]
  wire [5:0] Funct6D = io1_InstrD[31:26]; // @[cu.scala 66:29]
  wire [5:0] immI_lo_lo_lo = {io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31]}
    ; // @[Cat.scala 31:58]
  wire [12:0] immI_lo_lo = {io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],
    io1_InstrD[31],immI_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [25:0] immI_lo = {io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],
    io1_InstrD[31],immI_lo_lo_lo,immI_lo_lo}; // @[Cat.scala 31:58]
  wire [51:0] _immI_T_53 = {io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],io1_InstrD[31],
    io1_InstrD[31],immI_lo_lo_lo,immI_lo_lo,immI_lo}; // @[Cat.scala 31:58]
  wire [63:0] immI = {_immI_T_53,io1_InstrD[31:20]}; // @[Cat.scala 31:58]
  wire [11:0] _immS_T_2 = {Funct7D,io1_InstrD[11:7]}; // @[Cat.scala 31:58]
  wire [5:0] immS_lo_lo_lo = {_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11]}; // @[Cat.scala 31:58]
  wire [12:0] immS_lo_lo = {_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],
    _immS_T_2[11],immS_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [25:0] immS_lo = {_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[
    11],immS_lo_lo_lo,immS_lo_lo}; // @[Cat.scala 31:58]
  wire [51:0] _immS_T_55 = {_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],_immS_T_2[11],
    _immS_T_2[11],immS_lo_lo_lo,immS_lo_lo,immS_lo}; // @[Cat.scala 31:58]
  wire [63:0] immS = {_immS_T_55,Funct7D,io1_InstrD[11:7]}; // @[Cat.scala 31:58]
  wire [31:0] _immU_T_1 = {io1_InstrD[31:12],12'h0}; // @[Cat.scala 31:58]
  wire [7:0] immU_lo_lo = {_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1
    [31],_immU_T_1[31]}; // @[Cat.scala 31:58]
  wire [15:0] immU_lo = {_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1[
    31],_immU_T_1[31],immU_lo_lo}; // @[Cat.scala 31:58]
  wire [31:0] _immU_T_34 = {_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],_immU_T_1[31],
    _immU_T_1[31],_immU_T_1[31],immU_lo_lo,immU_lo}; // @[Cat.scala 31:58]
  wire [63:0] immU = {_immU_T_34,io1_InstrD[31:12],12'h0}; // @[Cat.scala 31:58]
  wire [12:0] _immSB_T_4 = {io1_InstrD[31],io1_InstrD[7],io1_InstrD[30:25],io1_InstrD[11:8],1'h0}; // @[Cat.scala 31:58]
  wire [5:0] immSB_lo_lo_lo = {_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12]
    }; // @[Cat.scala 31:58]
  wire [11:0] immSB_lo_lo = {_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],
    immSB_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [12:0] immSB_lo_hi = {_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],
    _immSB_T_4[12],immSB_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [24:0] immSB_lo_1 = {_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],
    _immSB_T_4[12],immSB_lo_lo_lo,immSB_lo_lo}; // @[Cat.scala 31:58]
  wire [50:0] _immSB_T_56 = {_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],
    _immSB_T_4[12],immSB_lo_lo_lo,immSB_lo_hi,immSB_lo_1}; // @[Cat.scala 31:58]
  wire [63:0] immSB = {_immSB_T_56,io1_InstrD[31],io1_InstrD[7],io1_InstrD[30:25],io1_InstrD[11:8],1'h0}; // @[Cat.scala 31:58]
  wire [19:0] immUJ = {io1_InstrD[31],io1_InstrD[19:12],io1_InstrD[20],io1_InstrD[30:21]}; // @[Cat.scala 31:58]
  wire [3:0] _inst_code_type_T_2 = 7'h0 == Funct7D ? 4'hf : 4'h0; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_4 = 6'h0 == Funct6D ? 5'h13 : 5'h0; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_6 = 6'h10 == Funct6D ? 5'h14 : _inst_code_type_T_4; // @[Mux.scala 81:58]
  wire [3:0] _inst_code_type_T_8 = 3'h2 == Funct3D ? 4'hd : 4'h4; // @[Mux.scala 81:58]
  wire [3:0] _inst_code_type_T_10 = 3'h3 == Funct3D ? 4'he : _inst_code_type_T_8; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_12 = 3'h4 == Funct3D ? 5'h17 : {{1'd0}, _inst_code_type_T_10}; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_14 = 3'h6 == Funct3D ? 5'h16 : _inst_code_type_T_12; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_16 = 3'h7 == Funct3D ? 5'h15 : _inst_code_type_T_14; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_18 = 3'h1 == Funct3D ? {{1'd0}, _inst_code_type_T_2} : _inst_code_type_T_16; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_20 = 3'h1 == Funct3D ? 5'hf : _inst_code_type_T_18; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_22 = 3'h5 == Funct3D ? _inst_code_type_T_6 : _inst_code_type_T_20; // @[Mux.scala 81:58]
  wire [7:0] _inst_code_type_T_23 = {_inst_code_type_T_22,3'h2}; // @[Cat.scala 31:58]
  wire [5:0] _inst_code_type_T_25 = 7'h20 == Funct7D ? 6'h36 : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_27 = 7'h0 == Funct7D ? 6'h30 : _inst_code_type_T_25; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_29 = 7'h1 == Funct7D ? 6'h2c : _inst_code_type_T_27; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_31 = 7'h0 == Funct7D ? 6'h31 : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_33 = 7'h1 == Funct7D ? 6'h2d : _inst_code_type_T_31; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_35 = 7'h1 == Funct7D ? 6'h2f : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_37 = 7'h0 == Funct7D ? 6'h34 : _inst_code_type_T_35; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_39 = 7'h0 == Funct7D ? 6'h35 : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_41 = 7'h1 == Funct7D ? 6'h2e : _inst_code_type_T_39; // @[Mux.scala 81:58]
  wire [6:0] _inst_code_type_T_43 = 7'h0 == Funct7D ? 7'h41 : 7'h0; // @[Mux.scala 81:58]
  wire [6:0] _inst_code_type_T_45 = 7'h1 == Funct7D ? 7'h24 : _inst_code_type_T_43; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_47 = 7'h0 == Funct7D ? 6'h32 : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_49 = 7'h1 == Funct7D ? 6'h23 : _inst_code_type_T_47; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_51 = 7'h20 == Funct7D ? 6'h33 : _inst_code_type_T_49; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_53 = 7'h0 == Funct7D ? 6'h38 : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_55 = 7'h1 == Funct7D ? 6'h26 : _inst_code_type_T_53; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_57 = 7'h0 == Funct7D ? 6'h37 : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_59 = 7'h1 == Funct7D ? 6'h25 : _inst_code_type_T_57; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_61 = 3'h1 == Funct3D ? _inst_code_type_T_33 : _inst_code_type_T_29; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_63 = 3'h2 == Funct3D ? _inst_code_type_T_37 : _inst_code_type_T_61; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_65 = 3'h3 == Funct3D ? _inst_code_type_T_41 : _inst_code_type_T_63; // @[Mux.scala 81:58]
  wire [6:0] _inst_code_type_T_67 = 3'h4 == Funct3D ? _inst_code_type_T_45 : {{1'd0}, _inst_code_type_T_65}; // @[Mux.scala 81:58]
  wire [6:0] _inst_code_type_T_69 = 3'h5 == Funct3D ? {{1'd0}, _inst_code_type_T_51} : _inst_code_type_T_67; // @[Mux.scala 81:58]
  wire [6:0] _inst_code_type_T_71 = 3'h6 == Funct3D ? {{1'd0}, _inst_code_type_T_55} : _inst_code_type_T_69; // @[Mux.scala 81:58]
  wire [6:0] _inst_code_type_T_73 = 3'h7 == Funct3D ? {{1'd0}, _inst_code_type_T_59} : _inst_code_type_T_71; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_74 = {_inst_code_type_T_73,3'h5}; // @[Cat.scala 31:58]
  wire [4:0] _inst_code_type_T_76 = 3'h0 == Funct3D ? 5'h1c : 5'h0; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_78 = 3'h1 == Funct3D ? 5'h1d : _inst_code_type_T_76; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_80 = 3'h4 == Funct3D ? 6'h20 : {{1'd0}, _inst_code_type_T_78}; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_82 = 3'h5 == Funct3D ? 6'h1e : _inst_code_type_T_80; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_84 = 3'h6 == Funct3D ? 6'h21 : _inst_code_type_T_82; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_86 = 3'h7 == Funct3D ? 6'h1f : _inst_code_type_T_84; // @[Mux.scala 81:58]
  wire [8:0] _inst_code_type_T_87 = {_inst_code_type_T_86,3'h4}; // @[Cat.scala 31:58]
  wire [3:0] _inst_code_type_T_93 = 3'h0 == Funct3D ? 4'h8 : 4'h0; // @[Mux.scala 81:58]
  wire [3:0] _inst_code_type_T_95 = 3'h1 == Funct3D ? 4'ha : _inst_code_type_T_93; // @[Mux.scala 81:58]
  wire [3:0] _inst_code_type_T_97 = 3'h2 == Funct3D ? 4'hc : _inst_code_type_T_95; // @[Mux.scala 81:58]
  wire [3:0] _inst_code_type_T_99 = 3'h4 == Funct3D ? 4'h7 : _inst_code_type_T_97; // @[Mux.scala 81:58]
  wire [3:0] _inst_code_type_T_101 = 3'h5 == Funct3D ? 4'h9 : _inst_code_type_T_99; // @[Mux.scala 81:58]
  wire [3:0] _inst_code_type_T_103 = 3'h6 == Funct3D ? 4'hb : _inst_code_type_T_101; // @[Mux.scala 81:58]
  wire [3:0] _inst_code_type_T_105 = 3'h3 == Funct3D ? 4'h6 : _inst_code_type_T_103; // @[Mux.scala 81:58]
  wire [6:0] _inst_code_type_T_106 = {_inst_code_type_T_105,3'h2}; // @[Cat.scala 31:58]
  wire [4:0] _inst_code_type_T_108 = 3'h0 == Funct3D ? 5'h18 : 5'h0; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_110 = 3'h1 == Funct3D ? 5'h19 : _inst_code_type_T_108; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_112 = 3'h2 == Funct3D ? 5'h1a : _inst_code_type_T_110; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_114 = 3'h3 == Funct3D ? 5'h1b : _inst_code_type_T_112; // @[Mux.scala 81:58]
  wire [7:0] _inst_code_type_T_115 = {_inst_code_type_T_114,3'h3}; // @[Cat.scala 31:58]
  wire [4:0] _inst_code_type_T_117 = 7'h0 == Funct7D ? 5'h11 : 5'h0; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_119 = 7'h20 == Funct7D ? 5'h12 : _inst_code_type_T_117; // @[Mux.scala 81:58]
  wire [2:0] _inst_code_type_T_121 = 3'h0 == Funct3D ? 3'h5 : 3'h0; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_123 = 3'h1 == Funct3D ? 5'h10 : {{2'd0}, _inst_code_type_T_121}; // @[Mux.scala 81:58]
  wire [4:0] _inst_code_type_T_125 = 3'h5 == Funct3D ? _inst_code_type_T_119 : _inst_code_type_T_123; // @[Mux.scala 81:58]
  wire [7:0] _inst_code_type_T_126 = {_inst_code_type_T_125,3'h2}; // @[Cat.scala 31:58]
  wire [5:0] _inst_code_type_T_128 = 7'h0 == Funct7D ? 6'h3c : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_130 = 7'h20 == Funct7D ? 6'h3d : _inst_code_type_T_128; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_132 = 7'h1 == Funct7D ? 6'h2b : _inst_code_type_T_130; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_134 = 7'h0 == Funct7D ? 6'h39 : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_136 = 7'h0 == Funct7D ? 6'h3a : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_138 = 7'h20 == Funct7D ? 6'h3b : _inst_code_type_T_136; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_140 = 7'h1 == Funct7D ? 6'h28 : _inst_code_type_T_138; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_142 = 3'h0 == Funct3D ? _inst_code_type_T_132 : 6'h0; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_144 = 3'h1 == Funct3D ? _inst_code_type_T_134 : _inst_code_type_T_142; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_146 = 3'h5 == Funct3D ? _inst_code_type_T_140 : _inst_code_type_T_144; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_148 = 3'h6 == Funct3D ? 6'h29 : _inst_code_type_T_146; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_150 = 3'h7 == Funct3D ? 6'h2a : _inst_code_type_T_148; // @[Mux.scala 81:58]
  wire [5:0] _inst_code_type_T_152 = 3'h4 == Funct3D ? 6'h27 : _inst_code_type_T_150; // @[Mux.scala 81:58]
  wire [8:0] _inst_code_type_T_153 = {_inst_code_type_T_152,3'h5}; // @[Cat.scala 31:58]
  wire [6:0] _inst_code_type_T_156 = 7'h0 == Funct7D ? 7'h4c : 7'h0; // @[Mux.scala 81:58]
  wire [6:0] _inst_code_type_T_158 = 7'h18 == Funct7D ? 7'h4d : _inst_code_type_T_156; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_159 = {_inst_code_type_T_158,3'h0}; // @[Cat.scala 31:58]
  wire [9:0] _inst_code_type_T_167 = 3'h0 == Funct3D ? _inst_code_type_T_159 : 10'h0; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_169 = 3'h1 == Funct3D ? 10'h25a : _inst_code_type_T_167; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_171 = 3'h2 == Funct3D ? 10'h252 : _inst_code_type_T_169; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_173 = 3'h3 == Funct3D ? 10'h24a : _inst_code_type_T_171; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_175 = 3'h5 == Funct3D ? 10'h242 : _inst_code_type_T_173; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_177 = 3'h6 == Funct3D ? 10'h23a : _inst_code_type_T_175; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_179 = 3'h7 == Funct3D ? 10'h232 : _inst_code_type_T_177; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_182 = 3'h1 == Funct3D ? 10'h277 : 10'h0; // @[Mux.scala 81:58]
  wire [7:0] _inst_code_type_T_184 = 7'h13 == OpD ? _inst_code_type_T_23 : 8'h0; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_186 = 7'h33 == OpD ? _inst_code_type_T_74 : {{2'd0}, _inst_code_type_T_184}; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_188 = 7'h63 == OpD ? {{1'd0}, _inst_code_type_T_87} : _inst_code_type_T_186; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_190 = 7'h6f == OpD ? 10'h16 : _inst_code_type_T_188; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_192 = 7'h67 == OpD ? 10'h1a : _inst_code_type_T_190; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_194 = 7'h37 == OpD ? 10'h9 : _inst_code_type_T_192; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_196 = 7'h17 == OpD ? 10'h201 : _inst_code_type_T_194; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_198 = 7'h3 == OpD ? {{3'd0}, _inst_code_type_T_106} : _inst_code_type_T_196; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_200 = 7'h23 == OpD ? {{2'd0}, _inst_code_type_T_115} : _inst_code_type_T_198; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_202 = 7'h1b == OpD ? {{2'd0}, _inst_code_type_T_126} : _inst_code_type_T_200; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_204 = 7'h3b == OpD ? {{1'd0}, _inst_code_type_T_153} : _inst_code_type_T_202; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_206 = 7'h0 == OpD ? 10'h282 : _inst_code_type_T_204; // @[Mux.scala 81:58]
  wire [9:0] _inst_code_type_T_208 = 7'h73 == OpD ? _inst_code_type_T_179 : _inst_code_type_T_206; // @[Mux.scala 81:58]
  wire [9:0] inst_code_type = 7'hf == OpD ? _inst_code_type_T_182 : _inst_code_type_T_208; // @[Mux.scala 81:58]
  wire [6:0] ins_code = inst_code_type[9:3]; // @[cu.scala 196:35]
  wire [2:0] inst_type = inst_code_type[2:0]; // @[cu.scala 197:35]
  wire [3:0] _io_csr_control_T_7 = 7'h4b == ins_code ? 4'h4 : 4'h0; // @[Mux.scala 81:58]
  wire [3:0] _io_csr_control_T_9 = 7'h48 == ins_code ? 4'h4 : _io_csr_control_T_7; // @[Mux.scala 81:58]
  wire [3:0] _io_csr_control_T_11 = 7'h49 == ins_code ? 4'h2 : _io_csr_control_T_9; // @[Mux.scala 81:58]
  wire [3:0] _io_csr_control_T_13 = 7'h46 == ins_code ? 4'h2 : _io_csr_control_T_11; // @[Mux.scala 81:58]
  wire [3:0] _io_csr_control_T_15 = 7'h4a == ins_code ? 4'h1 : _io_csr_control_T_13; // @[Mux.scala 81:58]
  wire [3:0] _io_csr_control_T_17 = 7'h47 == ins_code ? 4'h1 : _io_csr_control_T_15; // @[Mux.scala 81:58]
  wire  _io_ImmD_T = inst_type == 3'h1; // @[cu.scala 235:20]
  wire  _io_ImmD_T_1 = inst_type == 3'h2; // @[cu.scala 236:20]
  wire  _io_ImmD_T_2 = inst_type == 3'h3; // @[cu.scala 237:20]
  wire  _io_ImmD_T_3 = inst_type == 3'h4; // @[cu.scala 238:20]
  wire  _io_ImmD_T_4 = inst_type == 3'h6; // @[cu.scala 239:20]
  wire [63:0] _io_ImmD_T_5 = _io_ImmD_T ? immU : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_ImmD_T_6 = _io_ImmD_T_1 ? immI : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_ImmD_T_7 = _io_ImmD_T_2 ? immS : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_ImmD_T_8 = _io_ImmD_T_3 ? immSB : 64'h0; // @[Mux.scala 27:73]
  wire [19:0] _io_ImmD_T_9 = _io_ImmD_T_4 ? immUJ : 20'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_ImmD_T_10 = _io_ImmD_T_5 | _io_ImmD_T_6; // @[Mux.scala 27:73]
  wire [63:0] _io_ImmD_T_11 = _io_ImmD_T_10 | _io_ImmD_T_7; // @[Mux.scala 27:73]
  wire [63:0] _io_ImmD_T_12 = _io_ImmD_T_11 | _io_ImmD_T_8; // @[Mux.scala 27:73]
  wire [63:0] _GEN_0 = {{44'd0}, _io_ImmD_T_9}; // @[Mux.scala 27:73]
  wire  _io_RegWriteD_T_29 = 7'h30 == ins_code | (7'h2b == ins_code | (7'h2f == ins_code | (7'h2e == ins_code | (7'h2d
     == ins_code | (7'h2c == ins_code | (7'h2b == ins_code | (7'h2a == ins_code | (7'h29 == ins_code | (7'h28 ==
    ins_code | (7'h27 == ins_code | (7'h26 == ins_code | (7'h25 == ins_code | (7'h24 == ins_code | 7'h23 == ins_code))))
    ))))))))); // @[Mux.scala 81:58]
  wire  _io_RegWriteD_T_59 = 7'h2 == ins_code | (7'h3 == ins_code | (7'h3d == ins_code | (7'h3c == ins_code | (7'h3b ==
    ins_code | (7'h3a == ins_code | (7'h39 == ins_code | (7'h38 == ins_code | (7'h37 == ins_code | (7'h36 == ins_code |
    (7'h35 == ins_code | (7'h34 == ins_code | (7'h33 == ins_code | (7'h32 == ins_code | (7'h31 == ins_code |
    _io_RegWriteD_T_29)))))))))))))); // @[Mux.scala 81:58]
  wire  _io_RegWriteD_T_89 = 7'h10 == ins_code | (7'hf == ins_code | (7'he == ins_code | (7'hd == ins_code | (7'h9 ==
    ins_code | (7'h7 == ins_code | (7'hc == ins_code | (7'hb == ins_code | (7'ha == ins_code | (7'h9 == ins_code | (7'h8
     == ins_code | (7'h7 == ins_code | (7'h6 == ins_code | (7'h5 == ins_code | (7'h4 == ins_code | _io_RegWriteD_T_59)))
    ))))))))))); // @[Mux.scala 81:58]
  wire  _io_RegWriteD_T_119 = 7'h47 == ins_code | (7'h48 == ins_code | (7'h4b == ins_code | (7'h4a == ins_code | (7'h49
     == ins_code | (7'h1 == ins_code | (7'h40 == ins_code | (7'h41 == ins_code | (7'h17 == ins_code | (7'h16 == ins_code
     | (7'h15 == ins_code | (7'h14 == ins_code | (7'h13 == ins_code | (7'h12 == ins_code | (7'h11 == ins_code |
    _io_RegWriteD_T_89)))))))))))))); // @[Mux.scala 81:58]
  wire  _io_ALUSrcD_1_T_4 = _io_ImmD_T_1 | _io_ImmD_T_4 | _io_ImmD_T; // @[cu.scala 363:79]
  wire [1:0] _io_ALUCtrlD_T_33 = 7'h40 == ins_code ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _io_ALUCtrlD_T_35 = 7'h30 == ins_code ? 2'h2 : _io_ALUCtrlD_T_33; // @[Mux.scala 81:58]
  wire [1:0] _io_ALUCtrlD_T_37 = 7'h5 == ins_code ? 2'h2 : _io_ALUCtrlD_T_35; // @[Mux.scala 81:58]
  wire [1:0] _io_ALUCtrlD_T_39 = 7'h4 == ins_code ? 2'h2 : _io_ALUCtrlD_T_37; // @[Mux.scala 81:58]
  wire [1:0] _io_ALUCtrlD_T_41 = 7'h3c == ins_code ? 2'h2 : _io_ALUCtrlD_T_39; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_43 = 7'hd == ins_code ? 16'h2000 : {{14'd0}, _io_ALUCtrlD_T_41}; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_45 = 7'he == ins_code ? 16'h4000 : _io_ALUCtrlD_T_43; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_47 = 7'hf == ins_code ? 16'h1000 : _io_ALUCtrlD_T_45; // @[Mux.scala 81:58]
  wire [15:0] _io_ALUCtrlD_T_49 = 7'h10 == ins_code ? 16'h1000 : _io_ALUCtrlD_T_47; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_51 = 7'h11 == ins_code ? 32'h10000 : {{16'd0}, _io_ALUCtrlD_T_49}; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_53 = 7'h12 == ins_code ? 32'h8000 : _io_ALUCtrlD_T_51; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_55 = 7'h13 == ins_code ? 32'h10000 : _io_ALUCtrlD_T_53; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_57 = 7'h14 == ins_code ? 32'h8000 : _io_ALUCtrlD_T_55; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_59 = 7'h15 == ins_code ? 32'h10 : _io_ALUCtrlD_T_57; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_61 = 7'h16 == ins_code ? 32'h800 : _io_ALUCtrlD_T_59; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_63 = 7'h17 == ins_code ? 32'h100000 : _io_ALUCtrlD_T_61; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_65 = 7'h1 == ins_code ? 32'h80 : _io_ALUCtrlD_T_63; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_67 = 7'h30 == ins_code ? 32'h2 : _io_ALUCtrlD_T_65; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_69 = 7'h31 == ins_code ? 32'h1000 : _io_ALUCtrlD_T_67; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_71 = 7'h32 == ins_code ? 32'h10000 : _io_ALUCtrlD_T_69; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_73 = 7'h33 == ins_code ? 32'h8000 : _io_ALUCtrlD_T_71; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_75 = 7'h34 == ins_code ? 32'h2000 : _io_ALUCtrlD_T_73; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_77 = 7'h35 == ins_code ? 32'h4000 : _io_ALUCtrlD_T_75; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_79 = 7'h36 == ins_code ? 32'h20000 : _io_ALUCtrlD_T_77; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_81 = 7'h37 == ins_code ? 32'h10 : _io_ALUCtrlD_T_79; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_83 = 7'h38 == ins_code ? 32'h800 : _io_ALUCtrlD_T_81; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_85 = 7'h39 == ins_code ? 32'h1000 : _io_ALUCtrlD_T_83; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_87 = 7'h3a == ins_code ? 32'h10000 : _io_ALUCtrlD_T_85; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_89 = 7'h3b == ins_code ? 32'h8000 : _io_ALUCtrlD_T_87; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_91 = 7'h3c == ins_code ? 32'h2 : _io_ALUCtrlD_T_89; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_93 = 7'h3d == ins_code ? 32'h20000 : _io_ALUCtrlD_T_91; // @[Mux.scala 81:58]
  wire [31:0] _io_ALUCtrlD_T_95 = 7'h41 == ins_code ? 32'h100000 : _io_ALUCtrlD_T_93; // @[Mux.scala 81:58]
  wire [1:0] _io_MemWidthD_T_5 = 3'h2 == Funct3D ? 2'h2 : {{1'd0}, 3'h1 == Funct3D}; // @[Mux.scala 81:58]
  wire [1:0] _io_MemWidthD_T_7 = 3'h4 == Funct3D ? 2'h0 : _io_MemWidthD_T_5; // @[Mux.scala 81:58]
  wire [1:0] _io_MemWidthD_T_9 = 3'h5 == Funct3D ? 2'h1 : _io_MemWidthD_T_7; // @[Mux.scala 81:58]
  wire [1:0] _io_MemWidthD_T_11 = 3'h6 == Funct3D ? 2'h2 : _io_MemWidthD_T_9; // @[Mux.scala 81:58]
  wire [1:0] _io_MemWidthD_T_13 = 3'h3 == Funct3D ? 2'h3 : _io_MemWidthD_T_11; // @[Mux.scala 81:58]
  wire [1:0] _io_MemWidthD_T_21 = 3'h3 == Funct3D ? 2'h3 : _io_MemWidthD_T_5; // @[Mux.scala 81:58]
  wire [1:0] _io_MemWidthD_T_23 = 7'h3 == OpD ? _io_MemWidthD_T_13 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _io_muldiv_control_T_14 = 7'h24 == ins_code ? 2'h2 : 2'h0; // @[Mux.scala 81:58]
  wire [1:0] _io_muldiv_control_T_16 = 7'h23 == ins_code ? 2'h1 : _io_muldiv_control_T_14; // @[Mux.scala 81:58]
  wire [3:0] _io_muldiv_control_T_18 = 7'h25 == ins_code ? 4'h4 : {{2'd0}, _io_muldiv_control_T_16}; // @[Mux.scala 81:58]
  wire [3:0] _io_muldiv_control_T_20 = 7'h26 == ins_code ? 4'h8 : _io_muldiv_control_T_18; // @[Mux.scala 81:58]
  wire [7:0] _io_muldiv_control_T_22 = 7'h27 == ins_code ? 8'h10 : {{4'd0}, _io_muldiv_control_T_20}; // @[Mux.scala 81:58]
  wire [7:0] _io_muldiv_control_T_24 = 7'h28 == ins_code ? 8'h20 : _io_muldiv_control_T_22; // @[Mux.scala 81:58]
  wire [7:0] _io_muldiv_control_T_26 = 7'h29 == ins_code ? 8'h40 : _io_muldiv_control_T_24; // @[Mux.scala 81:58]
  wire [7:0] _io_muldiv_control_T_28 = 7'h2a == ins_code ? 8'h80 : _io_muldiv_control_T_26; // @[Mux.scala 81:58]
  wire [15:0] _io_muldiv_control_T_30 = 7'h2b == ins_code ? 16'h100 : {{8'd0}, _io_muldiv_control_T_28}; // @[Mux.scala 81:58]
  wire [15:0] _io_muldiv_control_T_32 = 7'h2c == ins_code ? 16'h200 : _io_muldiv_control_T_30; // @[Mux.scala 81:58]
  wire [15:0] _io_muldiv_control_T_34 = 7'h2d == ins_code ? 16'h400 : _io_muldiv_control_T_32; // @[Mux.scala 81:58]
  wire [15:0] _io_muldiv_control_T_36 = 7'h2f == ins_code ? 16'h1000 : _io_muldiv_control_T_34; // @[Mux.scala 81:58]
  wire [15:0] _io_muldiv_control_T_38 = 7'h2e == ins_code ? 16'h800 : _io_muldiv_control_T_36; // @[Mux.scala 81:58]
  assign io1_BadInstrD = ins_code == 7'h0; // @[cu.scala 259:31]
  assign io1_SysCallD = ins_code == 7'h4c; // @[cu.scala 260:31]
  assign io1_EretD = ins_code == 7'h4d; // @[cu.scala 261:31]
  assign io1_dmem_addr_cal = 7'h23 == OpD ? 3'h3 == Funct3D | (3'h2 == Funct3D | (3'h1 == Funct3D | 3'h0 == Funct3D)) : 7'h3
     == OpD & (3'h3 == Funct3D | (3'h6 == Funct3D | (3'h5 == Funct3D | (3'h4 == Funct3D | (3'h2 == Funct3D | (3'h1 ==
    Funct3D | 3'h0 == Funct3D)))))); // @[Mux.scala 81:58]
  assign io_RegWriteD = 7'h46 == ins_code | _io_RegWriteD_T_119; // @[Mux.scala 81:58]
  assign io_MemToRegD = 7'h3 == OpD & (3'h3 == Funct3D | (3'h6 == Funct3D | (3'h5 == Funct3D | (3'h4 == Funct3D | (3'h2
     == Funct3D | (3'h1 == Funct3D | 3'h0 == Funct3D)))))); // @[Mux.scala 81:58]
  assign io_MemWriteD = 7'h23 == OpD & (3'h3 == Funct3D | (3'h2 == Funct3D | (3'h1 == Funct3D | 3'h0 == Funct3D))); // @[Mux.scala 81:58]
  assign io_ALUCtrlD = _io_ALUCtrlD_T_95[23:0]; // @[cu.scala 384:17]
  assign io_ALUSrcD_0 = {{1'd0}, ins_code == 7'h40}; // @[cu.scala 361:19]
  assign io_ALUSrcD_1 = {{1'd0}, _io_ALUSrcD_1_T_4}; // @[cu.scala 363:19]
  assign io_RegDstD = io1_InstrD[11:7]; // @[cu.scala 76:29]
  assign io_LinkD = ins_code == 7'h3 | ins_code == 7'h2; // @[cu.scala 241:38]
  assign io_csrWriteD = 7'h46 == ins_code | (7'h47 == ins_code | (7'h48 == ins_code | (7'h4b == ins_code | (7'h4a ==
    ins_code | 7'h49 == ins_code)))); // @[Mux.scala 81:58]
  assign io_csrToRegD = 7'h46 == ins_code | (7'h47 == ins_code | (7'h48 == ins_code | (7'h4b == ins_code | (7'h4a ==
    ins_code | 7'h49 == ins_code)))); // @[Mux.scala 81:58]
  assign io_LoadUnsignedD = 7'h3 == OpD & (3'h6 == Funct3D | (3'h5 == Funct3D | 3'h4 == Funct3D)); // @[Mux.scala 81:58]
  assign io_MemWidthD = 7'h23 == OpD ? _io_MemWidthD_T_21 : _io_MemWidthD_T_23; // @[Mux.scala 81:58]
  assign io_ImmD = _io_ImmD_T_12 | _GEN_0; // @[Mux.scala 27:73]
  assign io_ebreakD = io1_InstrD == 32'h100073; // @[cu.scala 262:33]
  assign io_data_wD = 7'h12 == ins_code | (7'h11 == ins_code | (7'h10 == ins_code | (7'h5 == ins_code | (7'h3d ==
    ins_code | (7'h3c == ins_code | (7'h3b == ins_code | (7'h3a == ins_code | (7'h39 == ins_code | (7'h2b == ins_code |
    (7'h2b == ins_code | (7'h2a == ins_code | (7'h29 == ins_code | (7'h28 == ins_code | 7'h27 == ins_code))))))))))))); // @[Mux.scala 81:58]
  assign io_muldiv_control = {{8'd0}, _io_muldiv_control_T_38}; // @[cu.scala 475:23]
  assign io_muldiv_cal = io_muldiv_control != 24'h0; // @[cu.scala 491:40]
  assign io_alu_cal = io_ALUCtrlD != 24'h0; // @[cu.scala 492:34]
  assign io_csr_control = {{2'd0}, _io_csr_control_T_17}; // @[cu.scala 216:20]
  assign io_csr_Imm = ins_code == 7'h48 | ins_code == 7'h46 | ins_code == 7'h47; // @[cu.scala 224:72]
  assign io_fence_i_control = io1_InstrD == 32'h100f; // @[cu.scala 199:39]
endmodule
module dmem(
  input         io_data_ok,
  input  [63:0] io_rdata,
  input  [63:0] io_Physisc_Address,
  input  [1:0]  io_WIDTH,
  input         io_SIGN,
  output [63:0] io_RD,
  output        io_data_pending
);
  wire [1:0] ra = io_Physisc_Address[1:0]; // @[dmem.scala 39:32]
  wire  third_ra = io_Physisc_Address[2]; // @[dmem.scala 40:38]
  wire [2:0] _io_RD_T_1 = {ra,io_SIGN}; // @[Cat.scala 31:58]
  wire [6:0] io_RD_lo_lo_lo = {io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39
    ]}; // @[Cat.scala 31:58]
  wire [13:0] io_RD_lo_lo = {io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],
    io_RD_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [27:0] io_RD_lo = {io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],
    io_RD_lo_lo_lo,io_RD_lo_lo}; // @[Cat.scala 31:58]
  wire [55:0] _io_RD_T_59 = {io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],io_rdata[39],
    io_RD_lo_lo_lo,io_RD_lo_lo,io_RD_lo}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_61 = {_io_RD_T_59,io_rdata[39:32]}; // @[Cat.scala 31:58]
  wire [8:0] _io_RD_T_64 = {1'h0,io_rdata[39:32]}; // @[Cat.scala 31:58]
  wire [6:0] io_RD_lo_lo_lo_1 = {io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[
    47]}; // @[Cat.scala 31:58]
  wire [13:0] io_RD_lo_lo_1 = {io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47
    ],io_RD_lo_lo_lo_1}; // @[Cat.scala 31:58]
  wire [27:0] io_RD_lo_1 = {io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],
    io_RD_lo_lo_lo_1,io_RD_lo_lo_1}; // @[Cat.scala 31:58]
  wire [55:0] _io_RD_T_122 = {io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47]
    ,io_RD_lo_lo_lo_1,io_RD_lo_lo_1,io_RD_lo_1}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_124 = {_io_RD_T_122,io_rdata[47:40]}; // @[Cat.scala 31:58]
  wire [8:0] _io_RD_T_127 = {1'h0,io_rdata[47:40]}; // @[Cat.scala 31:58]
  wire [6:0] io_RD_lo_lo_lo_2 = {io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[
    55]}; // @[Cat.scala 31:58]
  wire [13:0] io_RD_lo_lo_2 = {io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55
    ],io_RD_lo_lo_lo_2}; // @[Cat.scala 31:58]
  wire [27:0] io_RD_lo_2 = {io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],
    io_RD_lo_lo_lo_2,io_RD_lo_lo_2}; // @[Cat.scala 31:58]
  wire [55:0] _io_RD_T_185 = {io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55],io_rdata[55]
    ,io_RD_lo_lo_lo_2,io_RD_lo_lo_2,io_RD_lo_2}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_187 = {_io_RD_T_185,io_rdata[55:48]}; // @[Cat.scala 31:58]
  wire [8:0] _io_RD_T_190 = {1'h0,io_rdata[55:48]}; // @[Cat.scala 31:58]
  wire [6:0] io_RD_lo_lo_lo_3 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[
    63]}; // @[Cat.scala 31:58]
  wire [13:0] io_RD_lo_lo_3 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63
    ],io_RD_lo_lo_lo_3}; // @[Cat.scala 31:58]
  wire [27:0] io_RD_lo_3 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],
    io_RD_lo_lo_lo_3,io_RD_lo_lo_3}; // @[Cat.scala 31:58]
  wire [55:0] _io_RD_T_248 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63]
    ,io_RD_lo_lo_lo_3,io_RD_lo_lo_3,io_RD_lo_3}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_250 = {_io_RD_T_248,io_rdata[63:56]}; // @[Cat.scala 31:58]
  wire [8:0] _io_RD_T_253 = {1'h0,io_rdata[63:56]}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_255 = 3'h0 == _io_RD_T_1 ? {{55'd0}, _io_RD_T_64} : _io_RD_T_61; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_257 = 3'h3 == _io_RD_T_1 ? _io_RD_T_124 : _io_RD_T_255; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_259 = 3'h2 == _io_RD_T_1 ? {{55'd0}, _io_RD_T_127} : _io_RD_T_257; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_261 = 3'h5 == _io_RD_T_1 ? _io_RD_T_187 : _io_RD_T_259; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_263 = 3'h4 == _io_RD_T_1 ? {{55'd0}, _io_RD_T_190} : _io_RD_T_261; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_265 = 3'h7 == _io_RD_T_1 ? _io_RD_T_250 : _io_RD_T_263; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_267 = 3'h6 == _io_RD_T_1 ? {{55'd0}, _io_RD_T_253} : _io_RD_T_265; // @[Mux.scala 81:58]
  wire [6:0] io_RD_lo_lo_lo_4 = {io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7]}; // @[Cat.scala 31:58]
  wire [13:0] io_RD_lo_lo_4 = {io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],
    io_RD_lo_lo_lo_4}; // @[Cat.scala 31:58]
  wire [27:0] io_RD_lo_4 = {io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],
    io_RD_lo_lo_lo_4,io_RD_lo_lo_4}; // @[Cat.scala 31:58]
  wire [55:0] _io_RD_T_327 = {io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],io_rdata[7],
    io_RD_lo_lo_lo_4,io_RD_lo_lo_4,io_RD_lo_4}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_329 = {_io_RD_T_327,io_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [8:0] _io_RD_T_332 = {1'h0,io_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [6:0] io_RD_lo_lo_lo_5 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[
    15]}; // @[Cat.scala 31:58]
  wire [13:0] io_RD_lo_lo_5 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15
    ],io_RD_lo_lo_lo_5}; // @[Cat.scala 31:58]
  wire [27:0] io_RD_lo_5 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],
    io_RD_lo_lo_lo_5,io_RD_lo_lo_5}; // @[Cat.scala 31:58]
  wire [55:0] _io_RD_T_390 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15]
    ,io_RD_lo_lo_lo_5,io_RD_lo_lo_5,io_RD_lo_5}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_392 = {_io_RD_T_390,io_rdata[15:8]}; // @[Cat.scala 31:58]
  wire [8:0] _io_RD_T_395 = {1'h0,io_rdata[15:8]}; // @[Cat.scala 31:58]
  wire [6:0] io_RD_lo_lo_lo_6 = {io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[
    23]}; // @[Cat.scala 31:58]
  wire [13:0] io_RD_lo_lo_6 = {io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23
    ],io_RD_lo_lo_lo_6}; // @[Cat.scala 31:58]
  wire [27:0] io_RD_lo_6 = {io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],
    io_RD_lo_lo_lo_6,io_RD_lo_lo_6}; // @[Cat.scala 31:58]
  wire [55:0] _io_RD_T_453 = {io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23],io_rdata[23]
    ,io_RD_lo_lo_lo_6,io_RD_lo_lo_6,io_RD_lo_6}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_455 = {_io_RD_T_453,io_rdata[23:16]}; // @[Cat.scala 31:58]
  wire [8:0] _io_RD_T_458 = {1'h0,io_rdata[23:16]}; // @[Cat.scala 31:58]
  wire [6:0] io_RD_lo_lo_lo_7 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[
    31]}; // @[Cat.scala 31:58]
  wire [13:0] io_RD_lo_lo_7 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31
    ],io_RD_lo_lo_lo_7}; // @[Cat.scala 31:58]
  wire [27:0] io_RD_lo_7 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],
    io_RD_lo_lo_lo_7,io_RD_lo_lo_7}; // @[Cat.scala 31:58]
  wire [55:0] _io_RD_T_516 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31]
    ,io_RD_lo_lo_lo_7,io_RD_lo_lo_7,io_RD_lo_7}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_518 = {_io_RD_T_516,io_rdata[31:24]}; // @[Cat.scala 31:58]
  wire [8:0] _io_RD_T_521 = {1'h0,io_rdata[31:24]}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_523 = 3'h0 == _io_RD_T_1 ? {{55'd0}, _io_RD_T_332} : _io_RD_T_329; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_525 = 3'h3 == _io_RD_T_1 ? _io_RD_T_392 : _io_RD_T_523; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_527 = 3'h2 == _io_RD_T_1 ? {{55'd0}, _io_RD_T_395} : _io_RD_T_525; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_529 = 3'h5 == _io_RD_T_1 ? _io_RD_T_455 : _io_RD_T_527; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_531 = 3'h4 == _io_RD_T_1 ? {{55'd0}, _io_RD_T_458} : _io_RD_T_529; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_533 = 3'h7 == _io_RD_T_1 ? _io_RD_T_518 : _io_RD_T_531; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_535 = 3'h6 == _io_RD_T_1 ? {{55'd0}, _io_RD_T_521} : _io_RD_T_533; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_536 = third_ra ? _io_RD_T_267 : _io_RD_T_535; // @[dmem.scala 72:19]
  wire [5:0] io_RD_lo_lo_lo_8 = {io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47]}; // @[Cat.scala 31:58]
  wire [11:0] io_RD_lo_lo_8 = {io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],
    io_RD_lo_lo_lo_8}; // @[Cat.scala 31:58]
  wire [23:0] io_RD_lo_8 = {io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],
    io_RD_lo_lo_lo_8,io_RD_lo_lo_8}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_590 = {io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],io_rdata[47],
    io_RD_lo_lo_lo_8,io_RD_lo_lo_8,io_RD_lo_8,io_rdata[47:32]}; // @[Cat.scala 31:58]
  wire [16:0] _io_RD_T_593 = {1'h0,io_rdata[47:32]}; // @[Cat.scala 31:58]
  wire [5:0] io_RD_lo_lo_lo_9 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63]}; // @[Cat.scala 31:58]
  wire [11:0] io_RD_lo_lo_9 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],
    io_RD_lo_lo_lo_9}; // @[Cat.scala 31:58]
  wire [23:0] io_RD_lo_9 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],
    io_RD_lo_lo_lo_9,io_RD_lo_lo_9}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_645 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],
    io_RD_lo_lo_lo_9,io_RD_lo_lo_9,io_RD_lo_9,io_rdata[63:48]}; // @[Cat.scala 31:58]
  wire [16:0] _io_RD_T_648 = {1'h0,io_rdata[63:48]}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_650 = 3'h1 == _io_RD_T_1 ? _io_RD_T_590 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_652 = 3'h0 == _io_RD_T_1 ? {{47'd0}, _io_RD_T_593} : _io_RD_T_650; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_654 = 3'h5 == _io_RD_T_1 ? _io_RD_T_645 : _io_RD_T_652; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_656 = 3'h4 == _io_RD_T_1 ? {{47'd0}, _io_RD_T_648} : _io_RD_T_654; // @[Mux.scala 81:58]
  wire [5:0] io_RD_lo_lo_lo_10 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15]}; // @[Cat.scala 31:58]
  wire [11:0] io_RD_lo_lo_10 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],
    io_RD_lo_lo_lo_10}; // @[Cat.scala 31:58]
  wire [23:0] io_RD_lo_10 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],
    io_RD_lo_lo_lo_10,io_RD_lo_lo_10}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_710 = {io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],io_rdata[15],
    io_RD_lo_lo_lo_10,io_RD_lo_lo_10,io_RD_lo_10,io_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [16:0] _io_RD_T_713 = {1'h0,io_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [5:0] io_RD_lo_lo_lo_11 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31]}; // @[Cat.scala 31:58]
  wire [11:0] io_RD_lo_lo_11 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],
    io_RD_lo_lo_lo_11}; // @[Cat.scala 31:58]
  wire [23:0] io_RD_lo_11 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],
    io_RD_lo_lo_lo_11,io_RD_lo_lo_11}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_765 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],
    io_RD_lo_lo_lo_11,io_RD_lo_lo_11,io_RD_lo_11,io_rdata[31:16]}; // @[Cat.scala 31:58]
  wire [16:0] _io_RD_T_768 = {1'h0,io_rdata[31:16]}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_770 = 3'h1 == _io_RD_T_1 ? _io_RD_T_710 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_772 = 3'h0 == _io_RD_T_1 ? {{47'd0}, _io_RD_T_713} : _io_RD_T_770; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_774 = 3'h5 == _io_RD_T_1 ? _io_RD_T_765 : _io_RD_T_772; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_776 = 3'h4 == _io_RD_T_1 ? {{47'd0}, _io_RD_T_768} : _io_RD_T_774; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_777 = third_ra ? _io_RD_T_656 : _io_RD_T_776; // @[dmem.scala 73:19]
  wire [7:0] io_RD_lo_lo_12 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63
    ],io_rdata[63]}; // @[Cat.scala 31:58]
  wire [15:0] io_RD_lo_12 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],
    io_rdata[63],io_RD_lo_lo_12}; // @[Cat.scala 31:58]
  wire [31:0] _io_RD_T_812 = {io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63],io_rdata[63]
    ,io_rdata[63],io_RD_lo_lo_12,io_RD_lo_12}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_814 = {_io_RD_T_812,io_rdata[63:32]}; // @[Cat.scala 31:58]
  wire [32:0] _io_RD_T_816 = {1'h0,io_rdata[63:32]}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_817 = io_SIGN ? _io_RD_T_814 : {{31'd0}, _io_RD_T_816}; // @[dmem.scala 65:12]
  wire [7:0] io_RD_lo_lo_13 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31
    ],io_rdata[31]}; // @[Cat.scala 31:58]
  wire [15:0] io_RD_lo_13 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],
    io_rdata[31],io_RD_lo_lo_13}; // @[Cat.scala 31:58]
  wire [31:0] _io_RD_T_852 = {io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31],io_rdata[31]
    ,io_rdata[31],io_RD_lo_lo_13,io_RD_lo_13}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_854 = {_io_RD_T_852,io_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [32:0] _io_RD_T_856 = {1'h0,io_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _io_RD_T_857 = io_SIGN ? _io_RD_T_854 : {{31'd0}, _io_RD_T_856}; // @[dmem.scala 65:12]
  wire [63:0] _io_RD_T_858 = third_ra ? _io_RD_T_817 : _io_RD_T_857; // @[dmem.scala 74:19]
  wire [63:0] _io_RD_T_860 = 2'h1 == io_WIDTH ? _io_RD_T_777 : _io_RD_T_536; // @[Mux.scala 81:58]
  wire [63:0] _io_RD_T_862 = 2'h2 == io_WIDTH ? _io_RD_T_858 : _io_RD_T_860; // @[Mux.scala 81:58]
  assign io_RD = 2'h3 == io_WIDTH ? io_rdata : _io_RD_T_862; // @[Mux.scala 81:58]
  assign io_data_pending = ~io_data_ok; // @[dmem.scala 36:24]
endmodule
module dmemreq(
  input         io_en,
  input         io_MemWriteE,
  input         io_MemToRegE,
  input  [1:0]  io_MemWidthE,
  input  [63:0] io_VAddrE,
  input  [63:0] io_WriteDataE,
  output        io_req,
  output        io_wr,
  output [1:0]  io_size,
  output [63:0] io_addr,
  output [63:0] io_wdata,
  output [7:0]  io_wstrb
);
  wire [2:0] ra = io_VAddrE[2:0]; // @[dmemreq.scala 99:23]
  wire [1:0] _io_wstrb_T_1 = 3'h1 == ra ? 2'h2 : 2'h1; // @[Mux.scala 81:58]
  wire [2:0] _io_wstrb_T_3 = 3'h2 == ra ? 3'h4 : {{1'd0}, _io_wstrb_T_1}; // @[Mux.scala 81:58]
  wire [3:0] _io_wstrb_T_5 = 3'h3 == ra ? 4'h8 : {{1'd0}, _io_wstrb_T_3}; // @[Mux.scala 81:58]
  wire [4:0] _io_wstrb_T_7 = 3'h4 == ra ? 5'h10 : {{1'd0}, _io_wstrb_T_5}; // @[Mux.scala 81:58]
  wire [5:0] _io_wstrb_T_9 = 3'h5 == ra ? 6'h20 : {{1'd0}, _io_wstrb_T_7}; // @[Mux.scala 81:58]
  wire [6:0] _io_wstrb_T_11 = 3'h6 == ra ? 7'h40 : {{1'd0}, _io_wstrb_T_9}; // @[Mux.scala 81:58]
  wire [7:0] _io_wstrb_T_13 = 3'h7 == ra ? 8'h80 : {{1'd0}, _io_wstrb_T_11}; // @[Mux.scala 81:58]
  wire [1:0] _io_wstrb_T_15 = 3'h0 == ra ? 2'h3 : 2'h0; // @[Mux.scala 81:58]
  wire [3:0] _io_wstrb_T_17 = 3'h2 == ra ? 4'hc : {{2'd0}, _io_wstrb_T_15}; // @[Mux.scala 81:58]
  wire [5:0] _io_wstrb_T_19 = 3'h4 == ra ? 6'h30 : {{2'd0}, _io_wstrb_T_17}; // @[Mux.scala 81:58]
  wire [7:0] _io_wstrb_T_21 = 3'h6 == ra ? 8'hc0 : {{2'd0}, _io_wstrb_T_19}; // @[Mux.scala 81:58]
  wire [3:0] _io_wstrb_T_23 = 3'h0 == ra ? 4'hf : 4'h0; // @[Mux.scala 81:58]
  wire [7:0] _io_wstrb_T_25 = 3'h4 == ra ? 8'hf0 : {{4'd0}, _io_wstrb_T_23}; // @[Mux.scala 81:58]
  wire [7:0] _io_wstrb_T_27 = 3'h0 == ra ? 8'hff : 8'h0; // @[Mux.scala 81:58]
  wire [7:0] _io_wstrb_T_29 = 2'h1 == io_MemWidthE ? _io_wstrb_T_21 : _io_wstrb_T_13; // @[Mux.scala 81:58]
  wire [7:0] _io_wstrb_T_31 = 2'h2 == io_MemWidthE ? _io_wstrb_T_25 : _io_wstrb_T_29; // @[Mux.scala 81:58]
  wire  _io_wdata_T_1 = io_VAddrE[31:29] == 3'h4; // @[macros.scala 479:55]
  wire [8:0] _io_wdata_T_5 = {1'h0,io_WriteDataE[7:0]}; // @[Cat.scala 31:58]
  wire [16:0] _io_wdata_T_9 = {1'h0,io_WriteDataE[7:0],8'h0}; // @[Cat.scala 31:58]
  wire [24:0] _io_wdata_T_13 = {1'h0,io_WriteDataE[7:0],16'h0}; // @[Cat.scala 31:58]
  wire [32:0] _io_wdata_T_17 = {1'h0,io_WriteDataE[7:0],24'h0}; // @[Cat.scala 31:58]
  wire [40:0] _io_wdata_T_21 = {1'h0,io_WriteDataE[7:0],32'h0}; // @[Cat.scala 31:58]
  wire [48:0] _io_wdata_T_25 = {1'h0,io_WriteDataE[7:0],40'h0}; // @[Cat.scala 31:58]
  wire [56:0] _io_wdata_T_29 = {1'h0,io_WriteDataE[7:0],48'h0}; // @[Cat.scala 31:58]
  wire [64:0] _io_wdata_T_33 = {1'h0,io_WriteDataE[7:0],56'h0}; // @[Cat.scala 31:58]
  wire [16:0] _io_wdata_T_35 = 3'h1 == ra ? _io_wdata_T_9 : {{8'd0}, _io_wdata_T_5}; // @[Mux.scala 81:58]
  wire [24:0] _io_wdata_T_37 = 3'h2 == ra ? _io_wdata_T_13 : {{8'd0}, _io_wdata_T_35}; // @[Mux.scala 81:58]
  wire [32:0] _io_wdata_T_39 = 3'h3 == ra ? _io_wdata_T_17 : {{8'd0}, _io_wdata_T_37}; // @[Mux.scala 81:58]
  wire [40:0] _io_wdata_T_41 = 3'h4 == ra ? _io_wdata_T_21 : {{8'd0}, _io_wdata_T_39}; // @[Mux.scala 81:58]
  wire [48:0] _io_wdata_T_43 = 3'h5 == ra ? _io_wdata_T_25 : {{8'd0}, _io_wdata_T_41}; // @[Mux.scala 81:58]
  wire [56:0] _io_wdata_T_45 = 3'h6 == ra ? _io_wdata_T_29 : {{8'd0}, _io_wdata_T_43}; // @[Mux.scala 81:58]
  wire [64:0] _io_wdata_T_47 = 3'h7 == ra ? _io_wdata_T_33 : {{8'd0}, _io_wdata_T_45}; // @[Mux.scala 81:58]
  wire [16:0] _io_wdata_T_50 = {1'h0,io_WriteDataE[15:0]}; // @[Cat.scala 31:58]
  wire [32:0] _io_wdata_T_54 = {1'h0,io_WriteDataE[15:0],16'h0}; // @[Cat.scala 31:58]
  wire [48:0] _io_wdata_T_58 = {1'h0,io_WriteDataE[15:0],32'h0}; // @[Cat.scala 31:58]
  wire [64:0] _io_wdata_T_62 = {1'h0,io_WriteDataE[15:0],48'h0}; // @[Cat.scala 31:58]
  wire [16:0] _io_wdata_T_64 = 3'h0 == ra ? _io_wdata_T_50 : 17'h0; // @[Mux.scala 81:58]
  wire [32:0] _io_wdata_T_66 = 3'h2 == ra ? _io_wdata_T_54 : {{16'd0}, _io_wdata_T_64}; // @[Mux.scala 81:58]
  wire [48:0] _io_wdata_T_68 = 3'h4 == ra ? _io_wdata_T_58 : {{16'd0}, _io_wdata_T_66}; // @[Mux.scala 81:58]
  wire [64:0] _io_wdata_T_70 = 3'h6 == ra ? _io_wdata_T_62 : {{16'd0}, _io_wdata_T_68}; // @[Mux.scala 81:58]
  wire [32:0] _io_wdata_T_73 = {1'h0,io_WriteDataE[31:0]}; // @[Cat.scala 31:58]
  wire [64:0] _io_wdata_T_77 = {1'h0,io_WriteDataE[31:0],32'h0}; // @[Cat.scala 31:58]
  wire [32:0] _io_wdata_T_79 = 3'h0 == ra ? _io_wdata_T_73 : 33'h0; // @[Mux.scala 81:58]
  wire [64:0] _io_wdata_T_81 = 3'h4 == ra ? _io_wdata_T_77 : {{32'd0}, _io_wdata_T_79}; // @[Mux.scala 81:58]
  wire [63:0] _io_wdata_T_83 = ra == 3'h0 ? io_WriteDataE : 64'h0; // @[dmemreq.scala 67:23]
  wire [64:0] _io_wdata_T_85 = 2'h1 == io_MemWidthE ? _io_wdata_T_70 : _io_wdata_T_47; // @[Mux.scala 81:58]
  wire [64:0] _io_wdata_T_87 = 2'h2 == io_MemWidthE ? _io_wdata_T_81 : _io_wdata_T_85; // @[Mux.scala 81:58]
  wire [64:0] _io_wdata_T_89 = 2'h3 == io_MemWidthE ? {{1'd0}, _io_wdata_T_83} : _io_wdata_T_87; // @[Mux.scala 81:58]
  wire [64:0] _io_wdata_T_90 = _io_wdata_T_1 ? _io_wdata_T_89 : {{1'd0}, io_WriteDataE}; // @[dmemreq.scala 114:23]
  assign io_req = io_en & (io_MemToRegE | io_MemWriteE); // @[dmemreq.scala 115:33]
  assign io_wr = io_MemWriteE; // @[dmemreq.scala 101:17]
  assign io_size = io_MemWidthE; // @[dmemreq.scala 111:17]
  assign io_addr = io_VAddrE; // @[dmemreq.scala 112:17]
  assign io_wdata = _io_wdata_T_90[63:0]; // @[dmemreq.scala 114:17]
  assign io_wstrb = 2'h3 == io_MemWidthE ? _io_wstrb_T_27 : _io_wstrb_T_31; // @[Mux.scala 81:58]
endmodule
module ex2mem(
  input         clock,
  input         reset,
  input         io1_RegWriteE,
  input         io1_MemToRegE,
  input         io1_LoadUnsignedE,
  input  [1:0]  io1_MemWidthE,
  input         io1_csrWriteE,
  input  [11:0] io1_WritecsrAddrE,
  input  [63:0] io1_PCE,
  input  [1:0]  io1_MemRLE,
  input  [1:0]  io1_BranchJump_JrE,
  input  [2:0]  io1_Tlb_Control,
  input         io1_eBreakE,
  input         io1_fence_i_control,
  input         io_en,
  input         io_clr,
  input  [63:0] io_WriteDataE,
  input  [4:0]  io_WriteRegE,
  input  [63:0] io_PhyAddrE,
  input  [63:0] io_CsrWritedataE,
  input  [31:0] io_ExceptionTypeE,
  input  [63:0] io_RtE,
  input  [63:0] io_Pc_NextE,
  input  [63:0] io_mem_trace_budleE_pc,
  input  [63:0] io_mem_trace_budleE_data,
  input  [1:0]  io_mem_trace_budleE_mem_fetch_type,
  input  [63:0] io_mem_trace_budleE_addr,
  input  [2:0]  io_mem_trace_budleE_len,
  input         io_mem_trace_budleE_cache,
  output        io_RegWriteM,
  output        io_MemToRegM,
  output [63:0] io_WriteDataM,
  output [4:0]  io_WriteRegM,
  output        io_LoadUnsignedM,
  output [1:0]  io_MemWidthM,
  output [63:0] io_PhyAddrM,
  output        io_csrWriteM,
  output [11:0] io_WritecsrAddrM,
  output [63:0] io_PCM,
  output [31:0] io_ExceptionTypeM_Out,
  output [1:0]  io_MemRLM,
  output [63:0] io_RtM,
  output [1:0]  io_BranchJump_JrM,
  output [2:0]  io_Tlb_ControlM,
  output        io_eBreakM,
  output [63:0] io_Pc_NextM,
  output [63:0] io_mem_trace_budleM_pc,
  output [63:0] io_mem_trace_budleM_data,
  output [1:0]  io_mem_trace_budleM_mem_fetch_type,
  output [63:0] io_mem_trace_budleM_addr,
  output [2:0]  io_mem_trace_budleM_len,
  output        io_mem_trace_budleM_cache,
  output [63:0] io_CsrWritedataM,
  output        io_fence_i_controlM
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [31:0] _RAND_24;
`endif // RANDOMIZE_REG_INIT
  reg  RegWrite_Reg; // @[ex2mem.scala 59:38]
  reg  MemToReg_Reg; // @[ex2mem.scala 60:38]
  reg [63:0] WriteData_Reg; // @[ex2mem.scala 63:39]
  reg [4:0] WriteReg_Reg; // @[ex2mem.scala 64:38]
  reg  LoadUnsigned_Reg; // @[ex2mem.scala 67:42]
  reg [1:0] MemWidth_Reg; // @[ex2mem.scala 68:38]
  reg [63:0] PhyAddr_Reg; // @[ex2mem.scala 69:37]
  reg  csrWrite_Reg; // @[ex2mem.scala 73:38]
  reg [11:0] WritecsrAddr_Reg; // @[ex2mem.scala 75:42]
  reg [63:0] PC_Reg; // @[ex2mem.scala 78:32]
  reg [31:0] ExceptionType_Reg; // @[ex2mem.scala 80:41]
  reg [1:0] MemRLM_Reg; // @[ex2mem.scala 81:40]
  reg [63:0] RtM_Reg; // @[ex2mem.scala 82:32]
  reg [1:0] BranchJump_JrM_Reg; // @[ex2mem.scala 83:43]
  reg [2:0] Tlb_Control_Reg; // @[ex2mem.scala 84:43]
  reg  eBreak_Reg; // @[ex2mem.scala 85:36]
  reg [63:0] pc_nextReg; // @[ex2mem.scala 86:36]
  reg [63:0] mem_trace_budleReg_pc; // @[ex2mem.scala 87:43]
  reg [63:0] mem_trace_budleReg_data; // @[ex2mem.scala 87:43]
  reg [1:0] mem_trace_budleReg_mem_fetch_type; // @[ex2mem.scala 87:43]
  reg [63:0] mem_trace_budleReg_addr; // @[ex2mem.scala 87:43]
  reg [2:0] mem_trace_budleReg_len; // @[ex2mem.scala 87:43]
  reg  mem_trace_budleReg_cache; // @[ex2mem.scala 87:43]
  reg [63:0] CsrWritedataReg; // @[ex2mem.scala 88:43]
  reg  fence_i_controlReg; // @[ex2mem.scala 90:43]
  assign io_RegWriteM = RegWrite_Reg; // @[ex2mem.scala 124:30]
  assign io_MemToRegM = MemToReg_Reg; // @[ex2mem.scala 125:30]
  assign io_WriteDataM = WriteData_Reg; // @[ex2mem.scala 128:30]
  assign io_WriteRegM = WriteReg_Reg; // @[ex2mem.scala 129:30]
  assign io_LoadUnsignedM = LoadUnsigned_Reg; // @[ex2mem.scala 132:30]
  assign io_MemWidthM = MemWidth_Reg; // @[ex2mem.scala 133:30]
  assign io_PhyAddrM = PhyAddr_Reg; // @[ex2mem.scala 134:30]
  assign io_csrWriteM = csrWrite_Reg; // @[ex2mem.scala 137:30]
  assign io_WritecsrAddrM = WritecsrAddr_Reg; // @[ex2mem.scala 139:30]
  assign io_PCM = PC_Reg; // @[ex2mem.scala 142:30]
  assign io_ExceptionTypeM_Out = ExceptionType_Reg; // @[ex2mem.scala 144:30]
  assign io_MemRLM = MemRLM_Reg; // @[ex2mem.scala 145:30]
  assign io_RtM = RtM_Reg; // @[ex2mem.scala 146:30]
  assign io_BranchJump_JrM = BranchJump_JrM_Reg; // @[ex2mem.scala 147:30]
  assign io_Tlb_ControlM = Tlb_Control_Reg; // @[ex2mem.scala 148:30]
  assign io_eBreakM = eBreak_Reg; // @[ex2mem.scala 149:30]
  assign io_Pc_NextM = pc_nextReg; // @[ex2mem.scala 150:30]
  assign io_mem_trace_budleM_pc = mem_trace_budleReg_pc; // @[ex2mem.scala 151:30]
  assign io_mem_trace_budleM_data = mem_trace_budleReg_data; // @[ex2mem.scala 151:30]
  assign io_mem_trace_budleM_mem_fetch_type = mem_trace_budleReg_mem_fetch_type; // @[ex2mem.scala 151:30]
  assign io_mem_trace_budleM_addr = mem_trace_budleReg_addr; // @[ex2mem.scala 151:30]
  assign io_mem_trace_budleM_len = mem_trace_budleReg_len; // @[ex2mem.scala 151:30]
  assign io_mem_trace_budleM_cache = mem_trace_budleReg_cache; // @[ex2mem.scala 151:30]
  assign io_CsrWritedataM = CsrWritedataReg; // @[ex2mem.scala 152:30]
  assign io_fence_i_controlM = fence_i_controlReg; // @[ex2mem.scala 153:30]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 93:38]
      RegWrite_Reg <= 1'h0;
    end else if (io_clr) begin // @[ex2mem.scala 93:61]
      RegWrite_Reg <= 1'h0;
    end else if (io_en) begin
      RegWrite_Reg <= io1_RegWriteE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 112:38]
      MemToReg_Reg <= 1'h0;
    end else if (io_clr) begin // @[ex2mem.scala 112:61]
      MemToReg_Reg <= 1'h0;
    end else if (io_en) begin
      MemToReg_Reg <= io1_MemToRegE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 96:38]
      WriteData_Reg <= 64'h0;
    end else if (io_clr) begin // @[ex2mem.scala 96:61]
      WriteData_Reg <= 64'h0;
    end else if (io_en) begin
      WriteData_Reg <= io_WriteDataE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 97:38]
      WriteReg_Reg <= 5'h0;
    end else if (io_clr) begin // @[ex2mem.scala 97:61]
      WriteReg_Reg <= 5'h0;
    end else if (io_en) begin
      WriteReg_Reg <= io_WriteRegE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 100:38]
      LoadUnsigned_Reg <= 1'h0;
    end else if (io_clr) begin // @[ex2mem.scala 100:61]
      LoadUnsigned_Reg <= 1'h0;
    end else if (io_en) begin
      LoadUnsigned_Reg <= io1_LoadUnsignedE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 101:38]
      MemWidth_Reg <= 2'h0;
    end else if (io_clr) begin // @[ex2mem.scala 101:61]
      MemWidth_Reg <= 2'h0;
    end else if (io_en) begin
      MemWidth_Reg <= io1_MemWidthE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 102:38]
      PhyAddr_Reg <= 64'h0;
    end else if (io_clr) begin // @[ex2mem.scala 102:61]
      PhyAddr_Reg <= 64'h0;
    end else if (io_en) begin
      PhyAddr_Reg <= io_PhyAddrE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 104:38]
      csrWrite_Reg <= 1'h0;
    end else if (io_clr) begin // @[ex2mem.scala 104:61]
      csrWrite_Reg <= 1'h0;
    end else if (io_en) begin
      csrWrite_Reg <= io1_csrWriteE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 106:38]
      WritecsrAddr_Reg <= 12'h0;
    end else if (io_clr) begin // @[ex2mem.scala 106:61]
      WritecsrAddr_Reg <= 12'h0;
    end else if (io_en) begin
      WritecsrAddr_Reg <= io1_WritecsrAddrE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 109:38]
      PC_Reg <= 64'h0;
    end else if (io_clr) begin // @[ex2mem.scala 109:61]
      PC_Reg <= 64'h0;
    end else if (io_en) begin
      PC_Reg <= io1_PCE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 111:38]
      ExceptionType_Reg <= 32'h0;
    end else if (io_clr) begin // @[ex2mem.scala 111:61]
      ExceptionType_Reg <= 32'h0;
    end else if (io_en) begin
      ExceptionType_Reg <= io_ExceptionTypeE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 113:38]
      MemRLM_Reg <= 2'h0;
    end else if (io_clr) begin // @[ex2mem.scala 113:61]
      MemRLM_Reg <= 2'h0;
    end else if (io_en) begin
      MemRLM_Reg <= io1_MemRLE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 114:38]
      RtM_Reg <= 64'h0;
    end else if (io_clr) begin // @[ex2mem.scala 114:60]
      RtM_Reg <= 64'h0;
    end else if (io_en) begin
      RtM_Reg <= io_RtE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 115:38]
      BranchJump_JrM_Reg <= 2'h0;
    end else if (io_clr) begin // @[ex2mem.scala 115:60]
      BranchJump_JrM_Reg <= 2'h0;
    end else if (io_en) begin
      BranchJump_JrM_Reg <= io1_BranchJump_JrE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 116:38]
      Tlb_Control_Reg <= 3'h0;
    end else if (io_clr) begin // @[ex2mem.scala 116:61]
      Tlb_Control_Reg <= 3'h0;
    end else if (io_en) begin
      Tlb_Control_Reg <= io1_Tlb_Control;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 117:38]
      eBreak_Reg <= 1'h0;
    end else if (io_clr) begin // @[ex2mem.scala 117:60]
      eBreak_Reg <= 1'h0;
    end else if (io_en) begin
      eBreak_Reg <= io1_eBreakE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 118:38]
      pc_nextReg <= 64'h0;
    end else if (io_clr) begin // @[ex2mem.scala 118:60]
      pc_nextReg <= 64'h0;
    end else if (io_en) begin
      pc_nextReg <= io_Pc_NextE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 119:38]
      mem_trace_budleReg_pc <= 64'h0;
    end else if (io_clr) begin // @[ex2mem.scala 119:97]
      mem_trace_budleReg_pc <= 64'h0;
    end else if (io_en) begin
      mem_trace_budleReg_pc <= io_mem_trace_budleE_pc;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 119:38]
      mem_trace_budleReg_data <= 64'h0;
    end else if (io_clr) begin // @[ex2mem.scala 119:97]
      mem_trace_budleReg_data <= 64'h0;
    end else if (io_en) begin
      mem_trace_budleReg_data <= io_mem_trace_budleE_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 119:38]
      mem_trace_budleReg_mem_fetch_type <= 2'h0;
    end else if (io_clr) begin // @[ex2mem.scala 119:97]
      mem_trace_budleReg_mem_fetch_type <= 2'h0;
    end else if (io_en) begin
      mem_trace_budleReg_mem_fetch_type <= io_mem_trace_budleE_mem_fetch_type;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 119:38]
      mem_trace_budleReg_addr <= 64'h0;
    end else if (io_clr) begin // @[ex2mem.scala 119:97]
      mem_trace_budleReg_addr <= 64'h0;
    end else if (io_en) begin
      mem_trace_budleReg_addr <= io_mem_trace_budleE_addr;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 119:38]
      mem_trace_budleReg_len <= 3'h0;
    end else if (io_clr) begin // @[ex2mem.scala 119:97]
      mem_trace_budleReg_len <= 3'h0;
    end else if (io_en) begin
      mem_trace_budleReg_len <= io_mem_trace_budleE_len;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 119:38]
      mem_trace_budleReg_cache <= 1'h0;
    end else if (io_clr) begin // @[ex2mem.scala 119:97]
      mem_trace_budleReg_cache <= 1'h0;
    end else if (io_en) begin
      mem_trace_budleReg_cache <= io_mem_trace_budleE_cache;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 120:38]
      CsrWritedataReg <= 64'h0;
    end else if (io_clr) begin // @[ex2mem.scala 120:60]
      CsrWritedataReg <= 64'h0;
    end else if (io_en) begin
      CsrWritedataReg <= io_CsrWritedataE;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ex2mem.scala 121:38]
      fence_i_controlReg <= 1'h0;
    end else if (io_clr) begin // @[ex2mem.scala 121:60]
      fence_i_controlReg <= 1'h0;
    end else if (io_en) begin
      fence_i_controlReg <= io1_fence_i_control;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  RegWrite_Reg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  MemToReg_Reg = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  WriteData_Reg = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  WriteReg_Reg = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  LoadUnsigned_Reg = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  MemWidth_Reg = _RAND_5[1:0];
  _RAND_6 = {2{`RANDOM}};
  PhyAddr_Reg = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  csrWrite_Reg = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  WritecsrAddr_Reg = _RAND_8[11:0];
  _RAND_9 = {2{`RANDOM}};
  PC_Reg = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  ExceptionType_Reg = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  MemRLM_Reg = _RAND_11[1:0];
  _RAND_12 = {2{`RANDOM}};
  RtM_Reg = _RAND_12[63:0];
  _RAND_13 = {1{`RANDOM}};
  BranchJump_JrM_Reg = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  Tlb_Control_Reg = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  eBreak_Reg = _RAND_15[0:0];
  _RAND_16 = {2{`RANDOM}};
  pc_nextReg = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  mem_trace_budleReg_pc = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  mem_trace_budleReg_data = _RAND_18[63:0];
  _RAND_19 = {1{`RANDOM}};
  mem_trace_budleReg_mem_fetch_type = _RAND_19[1:0];
  _RAND_20 = {2{`RANDOM}};
  mem_trace_budleReg_addr = _RAND_20[63:0];
  _RAND_21 = {1{`RANDOM}};
  mem_trace_budleReg_len = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  mem_trace_budleReg_cache = _RAND_22[0:0];
  _RAND_23 = {2{`RANDOM}};
  CsrWritedataReg = _RAND_23[63:0];
  _RAND_24 = {1{`RANDOM}};
  fence_i_controlReg = _RAND_24[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    RegWrite_Reg = 1'h0;
  end
  if (reset) begin
    MemToReg_Reg = 1'h0;
  end
  if (reset) begin
    WriteData_Reg = 64'h0;
  end
  if (reset) begin
    WriteReg_Reg = 5'h0;
  end
  if (reset) begin
    LoadUnsigned_Reg = 1'h0;
  end
  if (reset) begin
    MemWidth_Reg = 2'h0;
  end
  if (reset) begin
    PhyAddr_Reg = 64'h0;
  end
  if (reset) begin
    csrWrite_Reg = 1'h0;
  end
  if (reset) begin
    WritecsrAddr_Reg = 12'h0;
  end
  if (reset) begin
    PC_Reg = 64'h0;
  end
  if (reset) begin
    ExceptionType_Reg = 32'h0;
  end
  if (reset) begin
    MemRLM_Reg = 2'h0;
  end
  if (reset) begin
    RtM_Reg = 64'h0;
  end
  if (reset) begin
    BranchJump_JrM_Reg = 2'h0;
  end
  if (reset) begin
    Tlb_Control_Reg = 3'h0;
  end
  if (reset) begin
    eBreak_Reg = 1'h0;
  end
  if (reset) begin
    pc_nextReg = 64'h0;
  end
  if (reset) begin
    mem_trace_budleReg_pc = 64'h0;
  end
  if (reset) begin
    mem_trace_budleReg_data = 64'h0;
  end
  if (reset) begin
    mem_trace_budleReg_mem_fetch_type = 2'h0;
  end
  if (reset) begin
    mem_trace_budleReg_addr = 64'h0;
  end
  if (reset) begin
    mem_trace_budleReg_len = 3'h0;
  end
  if (reset) begin
    mem_trace_budleReg_cache = 1'h0;
  end
  if (reset) begin
    CsrWritedataReg = 64'h0;
  end
  if (reset) begin
    fence_i_controlReg = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module id2ex(
  input         clock,
  input         reset,
  input         io1_RegWriteD,
  input         io1_MemToRegD,
  input         io1_MemWriteD,
  input  [23:0] io1_ALUCtrlD,
  input  [1:0]  io1_ALUSrcD_0,
  input  [1:0]  io1_ALUSrcD_1,
  input  [4:0]  io1_RegDstD,
  input         io1_LinkD,
  input         io1_csrWriteD,
  input         io1_csrToRegD,
  input         io1_LoadUnsignedD,
  input  [1:0]  io1_MemWidthD,
  input         io1_ebreakD,
  input         io1_data_wD,
  input  [23:0] io1_muldiv_control,
  input         io1_muldiv_cal,
  input         io1_alu_cal,
  input  [5:0]  io1_csr_control,
  input         io1_csr_Imm,
  input         io1_fence_i_control,
  output        io2_RegWriteE,
  output        io2_MemToRegE,
  output        io2_MemWriteE,
  output [23:0] io2_ALUCtrlE,
  output        io2_ALUSrcE_0,
  output        io2_ALUSrcE_1,
  output [4:0]  io2_RegDstE,
  output        io2_LinkE,
  output [63:0] io2_PCPlus4E,
  output        io2_LoadUnsignedE,
  output [1:0]  io2_MemWidthE,
  output        io2_csrWriteE,
  output [11:0] io2_WritecsrAddrE,
  output [11:0] io2_ReadcsrAddrE,
  output [63:0] io2_PCE,
  output [1:0]  io2_BranchJump_JrE,
  output        io2_eBreakE,
  output        io2_fence_i_control,
  input         io_en,
  input         io_clr,
  output        io_csrToRegE_Out,
  input  [63:0] io_RD1D,
  input  [63:0] io_RD2D,
  input  [4:0]  io_R2D,
  input  [4:0]  io_R1D,
  input  [63:0] io_ImmD,
  input  [63:0] io_PCPlus4D,
  input  [11:0] io_WritecsrAddrD,
  input  [11:0] io_ReadcsrAddrD,
  input  [63:0] io_PCD,
  input  [31:0] io_ExceptionTypeD,
  input  [63:0] io_Pc_NextD,
  input  [1:0]  io_BranchJump_JrD,
  output [63:0] io_RD1E,
  output [63:0] io_RD2E,
  output [4:0]  io_R2E,
  output [4:0]  io_R1E,
  output [63:0] io_ImmE,
  output        io_data_wE,
  output [63:0] io_Pc_NextE,
  output [23:0] io_muldiv_control,
  output        io_alu_calE,
  output        io_muldiv_calE,
  output [31:0] io_ExceptionTypeE_Out,
  output [5:0]  io_csr_controlE,
  output        io_csr_ImmE
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] RD1E_Reg; // @[id2ex.scala 97:30]
  reg [63:0] RD2E_Reg; // @[id2ex.scala 98:30]
  reg [4:0] R2E_Reg; // @[id2ex.scala 99:29]
  reg [4:0] R1E_Reg; // @[id2ex.scala 100:29]
  reg [63:0] ImmE_Reg; // @[id2ex.scala 102:30]
  reg [63:0] PCPlus4E_Reg; // @[id2ex.scala 104:34]
  reg [11:0] WritecsrAddrE_Reg; // @[id2ex.scala 109:39]
  reg [11:0] ReadcsrAddrE_Reg; // @[id2ex.scala 110:38]
  reg [63:0] PCE_Reg; // @[id2ex.scala 111:29]
  reg [31:0] ExceptionTypeE_Reg; // @[id2ex.scala 112:40]
  reg [1:0] BranchJump_JrE_Reg; // @[id2ex.scala 114:40]
  reg [63:0] Pc_NextReg; // @[id2ex.scala 119:32]
  reg  decoder_port_reg_RegWriteD; // @[id2ex.scala 123:38]
  reg  decoder_port_reg_MemToRegD; // @[id2ex.scala 123:38]
  reg  decoder_port_reg_MemWriteD; // @[id2ex.scala 123:38]
  reg [23:0] decoder_port_reg_ALUCtrlD; // @[id2ex.scala 123:38]
  reg [1:0] decoder_port_reg_ALUSrcD_0; // @[id2ex.scala 123:38]
  reg [1:0] decoder_port_reg_ALUSrcD_1; // @[id2ex.scala 123:38]
  reg [4:0] decoder_port_reg_RegDstD; // @[id2ex.scala 123:38]
  reg  decoder_port_reg_LinkD; // @[id2ex.scala 123:38]
  reg  decoder_port_reg_csrWriteD; // @[id2ex.scala 123:38]
  reg  decoder_port_reg_csrToRegD; // @[id2ex.scala 123:38]
  reg  decoder_port_reg_LoadUnsignedD; // @[id2ex.scala 123:38]
  reg [1:0] decoder_port_reg_MemWidthD; // @[id2ex.scala 123:38]
  reg  decoder_port_reg_ebreakD; // @[id2ex.scala 123:38]
  reg  decoder_port_reg_data_wD; // @[id2ex.scala 123:38]
  reg [23:0] decoder_port_reg_muldiv_control; // @[id2ex.scala 123:38]
  reg  decoder_port_reg_muldiv_cal; // @[id2ex.scala 123:38]
  reg  decoder_port_reg_alu_cal; // @[id2ex.scala 123:38]
  reg [5:0] decoder_port_reg_csr_control; // @[id2ex.scala 123:38]
  reg  decoder_port_reg_csr_Imm; // @[id2ex.scala 123:38]
  reg  decoder_port_reg_fence_i_control; // @[id2ex.scala 123:38]
  assign io2_RegWriteE = decoder_port_reg_RegWriteD; // @[id2ex.scala 147:23]
  assign io2_MemToRegE = decoder_port_reg_MemToRegD; // @[id2ex.scala 148:23]
  assign io2_MemWriteE = decoder_port_reg_MemWriteD; // @[id2ex.scala 149:23]
  assign io2_ALUCtrlE = decoder_port_reg_ALUCtrlD; // @[id2ex.scala 150:23]
  assign io2_ALUSrcE_0 = decoder_port_reg_ALUSrcD_0[0]; // @[id2ex.scala 151:23]
  assign io2_ALUSrcE_1 = decoder_port_reg_ALUSrcD_1[0]; // @[id2ex.scala 151:23]
  assign io2_RegDstE = decoder_port_reg_RegDstD; // @[id2ex.scala 152:23]
  assign io2_LinkE = decoder_port_reg_LinkD; // @[id2ex.scala 159:23]
  assign io2_PCPlus4E = PCPlus4E_Reg; // @[id2ex.scala 160:23]
  assign io2_LoadUnsignedE = decoder_port_reg_LoadUnsignedD; // @[id2ex.scala 161:23]
  assign io2_MemWidthE = decoder_port_reg_MemWidthD; // @[id2ex.scala 162:23]
  assign io2_csrWriteE = decoder_port_reg_csrWriteD; // @[id2ex.scala 163:23]
  assign io2_WritecsrAddrE = WritecsrAddrE_Reg; // @[id2ex.scala 165:23]
  assign io2_ReadcsrAddrE = ReadcsrAddrE_Reg; // @[id2ex.scala 166:23]
  assign io2_PCE = PCE_Reg; // @[id2ex.scala 167:23]
  assign io2_BranchJump_JrE = BranchJump_JrE_Reg; // @[id2ex.scala 170:24]
  assign io2_eBreakE = decoder_port_reg_ebreakD; // @[id2ex.scala 174:23]
  assign io2_fence_i_control = decoder_port_reg_fence_i_control; // @[id2ex.scala 175:25]
  assign io_csrToRegE_Out = decoder_port_reg_csrToRegD; // @[id2ex.scala 164:26]
  assign io_RD1E = RD1E_Reg; // @[id2ex.scala 153:23]
  assign io_RD2E = RD2E_Reg; // @[id2ex.scala 154:23]
  assign io_R2E = R2E_Reg; // @[id2ex.scala 155:23]
  assign io_R1E = R1E_Reg; // @[id2ex.scala 156:23]
  assign io_ImmE = ImmE_Reg; // @[id2ex.scala 158:23]
  assign io_data_wE = decoder_port_reg_data_wD; // @[id2ex.scala 173:23]
  assign io_Pc_NextE = Pc_NextReg; // @[id2ex.scala 176:23]
  assign io_muldiv_control = decoder_port_reg_muldiv_control; // @[id2ex.scala 177:23]
  assign io_alu_calE = decoder_port_reg_alu_cal; // @[id2ex.scala 146:23]
  assign io_muldiv_calE = decoder_port_reg_muldiv_cal; // @[id2ex.scala 145:23]
  assign io_ExceptionTypeE_Out = ExceptionTypeE_Reg; // @[id2ex.scala 169:26]
  assign io_csr_controlE = decoder_port_reg_csr_control; // @[id2ex.scala 179:23]
  assign io_csr_ImmE = decoder_port_reg_csr_Imm; // @[id2ex.scala 180:23]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 126:42]
      RD1E_Reg <= 64'h0;
    end else if (io_clr) begin // @[id2ex.scala 126:64]
      RD1E_Reg <= 64'h0;
    end else if (io_en) begin
      RD1E_Reg <= io_RD1D;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 127:42]
      RD2E_Reg <= 64'h0;
    end else if (io_clr) begin // @[id2ex.scala 127:64]
      RD2E_Reg <= 64'h0;
    end else if (io_en) begin
      RD2E_Reg <= io_RD2D;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 128:42]
      R2E_Reg <= 5'h0;
    end else if (io_clr) begin // @[id2ex.scala 128:64]
      R2E_Reg <= 5'h0;
    end else if (io_en) begin
      R2E_Reg <= io_R2D;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 129:42]
      R1E_Reg <= 5'h0;
    end else if (io_clr) begin // @[id2ex.scala 129:64]
      R1E_Reg <= 5'h0;
    end else if (io_en) begin
      R1E_Reg <= io_R1D;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 131:42]
      ImmE_Reg <= 64'h0;
    end else if (io_clr) begin // @[id2ex.scala 131:64]
      ImmE_Reg <= 64'h0;
    end else if (io_en) begin
      ImmE_Reg <= io_ImmD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 132:42]
      PCPlus4E_Reg <= 64'h0;
    end else if (io_clr) begin // @[id2ex.scala 132:64]
      PCPlus4E_Reg <= 64'h0;
    end else if (io_en) begin
      PCPlus4E_Reg <= io_PCPlus4D;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 133:42]
      WritecsrAddrE_Reg <= 12'h0;
    end else if (io_clr) begin // @[id2ex.scala 133:64]
      WritecsrAddrE_Reg <= 12'h0;
    end else if (io_en) begin
      WritecsrAddrE_Reg <= io_WritecsrAddrD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 135:42]
      ReadcsrAddrE_Reg <= 12'h0;
    end else if (io_clr) begin // @[id2ex.scala 135:64]
      ReadcsrAddrE_Reg <= 12'h0;
    end else if (io_en) begin
      ReadcsrAddrE_Reg <= io_ReadcsrAddrD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 137:42]
      PCE_Reg <= 64'h0;
    end else if (io_clr) begin // @[id2ex.scala 137:64]
      PCE_Reg <= 64'h0;
    end else if (io_en) begin
      PCE_Reg <= io_PCD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 138:42]
      ExceptionTypeE_Reg <= 32'h0;
    end else if (io_clr) begin // @[id2ex.scala 138:64]
      ExceptionTypeE_Reg <= 32'h0;
    end else if (io_en) begin
      ExceptionTypeE_Reg <= io_ExceptionTypeD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 139:42]
      BranchJump_JrE_Reg <= 2'h0;
    end else if (io_clr) begin // @[id2ex.scala 139:64]
      BranchJump_JrE_Reg <= 2'h0;
    end else if (io_en) begin
      BranchJump_JrE_Reg <= io_BranchJump_JrD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 142:42]
      Pc_NextReg <= 64'h0;
    end else if (io_clr) begin // @[id2ex.scala 142:64]
      Pc_NextReg <= 64'h0;
    end else if (io_en) begin
      Pc_NextReg <= io_Pc_NextD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 124:28]
      decoder_port_reg_RegWriteD <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 124:77]
      decoder_port_reg_RegWriteD <= 1'h0;
    end else if (io_en) begin
      decoder_port_reg_RegWriteD <= io1_RegWriteD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 124:28]
      decoder_port_reg_MemToRegD <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 124:77]
      decoder_port_reg_MemToRegD <= 1'h0;
    end else if (io_en) begin
      decoder_port_reg_MemToRegD <= io1_MemToRegD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 124:28]
      decoder_port_reg_MemWriteD <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 124:77]
      decoder_port_reg_MemWriteD <= 1'h0;
    end else if (io_en) begin
      decoder_port_reg_MemWriteD <= io1_MemWriteD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 124:28]
      decoder_port_reg_ALUCtrlD <= 24'h0;
    end else if (io_clr) begin // @[id2ex.scala 124:77]
      decoder_port_reg_ALUCtrlD <= 24'h0;
    end else if (io_en) begin
      decoder_port_reg_ALUCtrlD <= io1_ALUCtrlD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 124:28]
      decoder_port_reg_ALUSrcD_0 <= 2'h0;
    end else if (io_clr) begin // @[id2ex.scala 124:77]
      decoder_port_reg_ALUSrcD_0 <= 2'h0;
    end else if (io_en) begin
      decoder_port_reg_ALUSrcD_0 <= io1_ALUSrcD_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 124:28]
      decoder_port_reg_ALUSrcD_1 <= 2'h0;
    end else if (io_clr) begin // @[id2ex.scala 124:77]
      decoder_port_reg_ALUSrcD_1 <= 2'h0;
    end else if (io_en) begin
      decoder_port_reg_ALUSrcD_1 <= io1_ALUSrcD_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 124:28]
      decoder_port_reg_RegDstD <= 5'h0;
    end else if (io_clr) begin // @[id2ex.scala 124:77]
      decoder_port_reg_RegDstD <= 5'h0;
    end else if (io_en) begin
      decoder_port_reg_RegDstD <= io1_RegDstD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 124:28]
      decoder_port_reg_LinkD <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 124:77]
      decoder_port_reg_LinkD <= 1'h0;
    end else if (io_en) begin
      decoder_port_reg_LinkD <= io1_LinkD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 124:28]
      decoder_port_reg_csrWriteD <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 124:77]
      decoder_port_reg_csrWriteD <= 1'h0;
    end else if (io_en) begin
      decoder_port_reg_csrWriteD <= io1_csrWriteD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 124:28]
      decoder_port_reg_csrToRegD <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 124:77]
      decoder_port_reg_csrToRegD <= 1'h0;
    end else if (io_en) begin
      decoder_port_reg_csrToRegD <= io1_csrToRegD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 124:28]
      decoder_port_reg_LoadUnsignedD <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 124:77]
      decoder_port_reg_LoadUnsignedD <= 1'h0;
    end else if (io_en) begin
      decoder_port_reg_LoadUnsignedD <= io1_LoadUnsignedD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 124:28]
      decoder_port_reg_MemWidthD <= 2'h0;
    end else if (io_clr) begin // @[id2ex.scala 124:77]
      decoder_port_reg_MemWidthD <= 2'h0;
    end else if (io_en) begin
      decoder_port_reg_MemWidthD <= io1_MemWidthD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 124:28]
      decoder_port_reg_ebreakD <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 124:77]
      decoder_port_reg_ebreakD <= 1'h0;
    end else if (io_en) begin
      decoder_port_reg_ebreakD <= io1_ebreakD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 124:28]
      decoder_port_reg_data_wD <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 124:77]
      decoder_port_reg_data_wD <= 1'h0;
    end else if (io_en) begin
      decoder_port_reg_data_wD <= io1_data_wD;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 124:28]
      decoder_port_reg_muldiv_control <= 24'h0;
    end else if (io_clr) begin // @[id2ex.scala 124:77]
      decoder_port_reg_muldiv_control <= 24'h0;
    end else if (io_en) begin
      decoder_port_reg_muldiv_control <= io1_muldiv_control;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 124:28]
      decoder_port_reg_muldiv_cal <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 124:77]
      decoder_port_reg_muldiv_cal <= 1'h0;
    end else if (io_en) begin
      decoder_port_reg_muldiv_cal <= io1_muldiv_cal;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 124:28]
      decoder_port_reg_alu_cal <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 124:77]
      decoder_port_reg_alu_cal <= 1'h0;
    end else if (io_en) begin
      decoder_port_reg_alu_cal <= io1_alu_cal;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 124:28]
      decoder_port_reg_csr_control <= 6'h0;
    end else if (io_clr) begin // @[id2ex.scala 124:77]
      decoder_port_reg_csr_control <= 6'h0;
    end else if (io_en) begin
      decoder_port_reg_csr_control <= io1_csr_control;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 124:28]
      decoder_port_reg_csr_Imm <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 124:77]
      decoder_port_reg_csr_Imm <= 1'h0;
    end else if (io_en) begin
      decoder_port_reg_csr_Imm <= io1_csr_Imm;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[id2ex.scala 124:28]
      decoder_port_reg_fence_i_control <= 1'h0;
    end else if (io_clr) begin // @[id2ex.scala 124:77]
      decoder_port_reg_fence_i_control <= 1'h0;
    end else if (io_en) begin
      decoder_port_reg_fence_i_control <= io1_fence_i_control;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  RD1E_Reg = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  RD2E_Reg = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  R2E_Reg = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  R1E_Reg = _RAND_3[4:0];
  _RAND_4 = {2{`RANDOM}};
  ImmE_Reg = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  PCPlus4E_Reg = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  WritecsrAddrE_Reg = _RAND_6[11:0];
  _RAND_7 = {1{`RANDOM}};
  ReadcsrAddrE_Reg = _RAND_7[11:0];
  _RAND_8 = {2{`RANDOM}};
  PCE_Reg = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  ExceptionTypeE_Reg = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  BranchJump_JrE_Reg = _RAND_10[1:0];
  _RAND_11 = {2{`RANDOM}};
  Pc_NextReg = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  decoder_port_reg_RegWriteD = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  decoder_port_reg_MemToRegD = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  decoder_port_reg_MemWriteD = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  decoder_port_reg_ALUCtrlD = _RAND_15[23:0];
  _RAND_16 = {1{`RANDOM}};
  decoder_port_reg_ALUSrcD_0 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  decoder_port_reg_ALUSrcD_1 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  decoder_port_reg_RegDstD = _RAND_18[4:0];
  _RAND_19 = {1{`RANDOM}};
  decoder_port_reg_LinkD = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  decoder_port_reg_csrWriteD = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  decoder_port_reg_csrToRegD = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  decoder_port_reg_LoadUnsignedD = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  decoder_port_reg_MemWidthD = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  decoder_port_reg_ebreakD = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  decoder_port_reg_data_wD = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  decoder_port_reg_muldiv_control = _RAND_26[23:0];
  _RAND_27 = {1{`RANDOM}};
  decoder_port_reg_muldiv_cal = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  decoder_port_reg_alu_cal = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  decoder_port_reg_csr_control = _RAND_29[5:0];
  _RAND_30 = {1{`RANDOM}};
  decoder_port_reg_csr_Imm = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  decoder_port_reg_fence_i_control = _RAND_31[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    RD1E_Reg = 64'h0;
  end
  if (reset) begin
    RD2E_Reg = 64'h0;
  end
  if (reset) begin
    R2E_Reg = 5'h0;
  end
  if (reset) begin
    R1E_Reg = 5'h0;
  end
  if (reset) begin
    ImmE_Reg = 64'h0;
  end
  if (reset) begin
    PCPlus4E_Reg = 64'h0;
  end
  if (reset) begin
    WritecsrAddrE_Reg = 12'h0;
  end
  if (reset) begin
    ReadcsrAddrE_Reg = 12'h0;
  end
  if (reset) begin
    PCE_Reg = 64'h0;
  end
  if (reset) begin
    ExceptionTypeE_Reg = 32'h0;
  end
  if (reset) begin
    BranchJump_JrE_Reg = 2'h0;
  end
  if (reset) begin
    Pc_NextReg = 64'h0;
  end
  if (reset) begin
    decoder_port_reg_RegWriteD = 1'h0;
  end
  if (reset) begin
    decoder_port_reg_MemToRegD = 1'h0;
  end
  if (reset) begin
    decoder_port_reg_MemWriteD = 1'h0;
  end
  if (reset) begin
    decoder_port_reg_ALUCtrlD = 24'h0;
  end
  if (reset) begin
    decoder_port_reg_ALUSrcD_0 = 2'h0;
  end
  if (reset) begin
    decoder_port_reg_ALUSrcD_1 = 2'h0;
  end
  if (reset) begin
    decoder_port_reg_RegDstD = 5'h0;
  end
  if (reset) begin
    decoder_port_reg_LinkD = 1'h0;
  end
  if (reset) begin
    decoder_port_reg_csrWriteD = 1'h0;
  end
  if (reset) begin
    decoder_port_reg_csrToRegD = 1'h0;
  end
  if (reset) begin
    decoder_port_reg_LoadUnsignedD = 1'h0;
  end
  if (reset) begin
    decoder_port_reg_MemWidthD = 2'h0;
  end
  if (reset) begin
    decoder_port_reg_ebreakD = 1'h0;
  end
  if (reset) begin
    decoder_port_reg_data_wD = 1'h0;
  end
  if (reset) begin
    decoder_port_reg_muldiv_control = 24'h0;
  end
  if (reset) begin
    decoder_port_reg_muldiv_cal = 1'h0;
  end
  if (reset) begin
    decoder_port_reg_alu_cal = 1'h0;
  end
  if (reset) begin
    decoder_port_reg_csr_control = 6'h0;
  end
  if (reset) begin
    decoder_port_reg_csr_Imm = 1'h0;
  end
  if (reset) begin
    decoder_port_reg_fence_i_control = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module if2id(
  input         clock,
  input         reset,
  input         io_en,
  input         io_clr,
  input  [63:0] io_InstrF,
  input  [63:0] io_PCPlus4F,
  input  [63:0] io_PCF,
  input  [1:0]  io_ExceptionTypeF,
  output [31:0] io_InstrD,
  output [63:0] io_PCPlus4D,
  output [63:0] io_PCD,
  output [1:0]  io_ExceptionTypeD_Out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] InstrD_Reg; // @[if2id.scala 30:29]
  reg [63:0] PCPlus4D_Reg; // @[if2id.scala 31:31]
  reg [63:0] PCD_Reg; // @[if2id.scala 33:26]
  reg [1:0] ExceptionTypeD_Reg; // @[if2id.scala 34:37]
  wire [63:0] _InstrD_Reg_T_2 = io_en ? io_InstrF : {{32'd0}, InstrD_Reg}; // @[if2id.scala 45:57]
  wire [63:0] _InstrD_Reg_T_3 = io_clr ? 64'h0 : _InstrD_Reg_T_2; // @[if2id.scala 45:35]
  assign io_InstrD = InstrD_Reg; // @[if2id.scala 38:15]
  assign io_PCPlus4D = PCPlus4D_Reg; // @[if2id.scala 39:17]
  assign io_PCD = PCD_Reg; // @[if2id.scala 42:13]
  assign io_ExceptionTypeD_Out = ExceptionTypeD_Reg; // @[if2id.scala 41:27]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[if2id.scala 30:29]
      InstrD_Reg <= 32'h13; // @[if2id.scala 30:29]
    end else begin
      InstrD_Reg <= _InstrD_Reg_T_3[31:0]; // @[if2id.scala 45:17]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[if2id.scala 46:35]
      PCPlus4D_Reg <= 64'h0;
    end else if (io_clr) begin // @[if2id.scala 46:57]
      PCPlus4D_Reg <= 64'h0;
    end else if (io_en) begin
      PCPlus4D_Reg <= io_PCPlus4F;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[if2id.scala 48:39]
      PCD_Reg <= 64'h0;
    end else if (io_clr) begin // @[if2id.scala 48:61]
      PCD_Reg <= 64'h0;
    end else if (io_en) begin
      PCD_Reg <= io_PCF;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[if2id.scala 49:39]
      ExceptionTypeD_Reg <= 2'h0;
    end else if (io_clr) begin // @[if2id.scala 49:61]
      ExceptionTypeD_Reg <= 2'h0;
    end else if (io_en) begin
      ExceptionTypeD_Reg <= io_ExceptionTypeF;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  InstrD_Reg = _RAND_0[31:0];
  _RAND_1 = {2{`RANDOM}};
  PCPlus4D_Reg = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  PCD_Reg = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  ExceptionTypeD_Reg = _RAND_3[1:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    InstrD_Reg = 32'h13;
  end
  if (reset) begin
    PCPlus4D_Reg = 64'h0;
  end
  if (reset) begin
    PCD_Reg = 64'h0;
  end
  if (reset) begin
    ExceptionTypeD_Reg = 2'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module mem2wb(
  input         clock,
  input         reset,
  input         io_en,
  input         io_clr,
  input         io_RegWriteM,
  input  [63:0] io_ResultM,
  input  [4:0]  io_WriteRegM,
  input         io_csrWriteM,
  input  [11:0] io_WritecsrAddrM,
  input  [63:0] io_CsrWritedataM,
  input  [63:0] io_PCM,
  input  [31:0] io_ExceptionTypeM,
  input  [1:0]  io_BranchJump_JrM,
  input         io_eBreakM,
  input  [63:0] io_Pc_NextM,
  input  [63:0] io_Mem_trace_budleM_pc,
  input  [63:0] io_Mem_trace_budleM_data,
  input  [1:0]  io_Mem_trace_budleM_mem_fetch_type,
  input  [63:0] io_Mem_trace_budleM_addr,
  input  [2:0]  io_Mem_trace_budleM_len,
  input         io_Mem_trace_budleM_cache,
  output        io_RegWriteW_Out,
  output [63:0] io_ResultW,
  output [4:0]  io_WriteRegW,
  output        io_csrWriteW,
  output [11:0] io_WritecsrAddrW,
  output [63:0] io_PCW,
  output [31:0] io_ExceptionTypeW_Out,
  output [1:0]  io_BranchJump_JrW,
  output        io_eBreakW,
  output [63:0] io_Pc_NextW,
  output [63:0] io_Mem_trace_budleW_pc,
  output [63:0] io_Mem_trace_budleW_data,
  output [1:0]  io_Mem_trace_budleW_mem_fetch_type,
  output [63:0] io_Mem_trace_budleW_addr,
  output [2:0]  io_Mem_trace_budleW_len,
  output        io_Mem_trace_budleW_cache,
  output [63:0] io_CsrWritedataW
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [63:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  reg  RegWriteW; // @[mem2wb.scala 51:34]
  reg [63:0] ResultW; // @[mem2wb.scala 54:32]
  reg [4:0] WriteRegW; // @[mem2wb.scala 55:34]
  reg  csrWriteW; // @[mem2wb.scala 57:34]
  reg [11:0] WritecsrAddrW; // @[mem2wb.scala 58:38]
  reg [63:0] PCW; // @[mem2wb.scala 60:28]
  reg [31:0] ExceptionTypeW; // @[mem2wb.scala 62:39]
  reg [1:0] BranchJump_JrW_Reg; // @[mem2wb.scala 64:43]
  reg  ebreak_Reg; // @[mem2wb.scala 66:40]
  reg [63:0] pc_nextReg; // @[mem2wb.scala 67:36]
  reg [63:0] Mem_trace_budleReg_pc; // @[mem2wb.scala 68:43]
  reg [63:0] Mem_trace_budleReg_data; // @[mem2wb.scala 68:43]
  reg [1:0] Mem_trace_budleReg_mem_fetch_type; // @[mem2wb.scala 68:43]
  reg [63:0] Mem_trace_budleReg_addr; // @[mem2wb.scala 68:43]
  reg [2:0] Mem_trace_budleReg_len; // @[mem2wb.scala 68:43]
  reg  Mem_trace_budleReg_cache; // @[mem2wb.scala 68:43]
  reg [63:0] CsrWritedataReg; // @[mem2wb.scala 69:40]
  assign io_RegWriteW_Out = RegWriteW; // @[mem2wb.scala 71:36]
  assign io_ResultW = ResultW; // @[mem2wb.scala 74:32]
  assign io_WriteRegW = WriteRegW; // @[mem2wb.scala 75:32]
  assign io_csrWriteW = csrWriteW; // @[mem2wb.scala 76:32]
  assign io_WritecsrAddrW = WritecsrAddrW; // @[mem2wb.scala 77:32]
  assign io_PCW = PCW; // @[mem2wb.scala 79:32]
  assign io_ExceptionTypeW_Out = ExceptionTypeW; // @[mem2wb.scala 81:32]
  assign io_BranchJump_JrW = BranchJump_JrW_Reg; // @[mem2wb.scala 82:32]
  assign io_eBreakW = ebreak_Reg; // @[mem2wb.scala 84:32]
  assign io_Pc_NextW = pc_nextReg; // @[mem2wb.scala 85:32]
  assign io_Mem_trace_budleW_pc = Mem_trace_budleReg_pc; // @[mem2wb.scala 86:33]
  assign io_Mem_trace_budleW_data = Mem_trace_budleReg_data; // @[mem2wb.scala 86:33]
  assign io_Mem_trace_budleW_mem_fetch_type = Mem_trace_budleReg_mem_fetch_type; // @[mem2wb.scala 86:33]
  assign io_Mem_trace_budleW_addr = Mem_trace_budleReg_addr; // @[mem2wb.scala 86:33]
  assign io_Mem_trace_budleW_len = Mem_trace_budleReg_len; // @[mem2wb.scala 86:33]
  assign io_Mem_trace_budleW_cache = Mem_trace_budleReg_cache; // @[mem2wb.scala 86:33]
  assign io_CsrWritedataW = CsrWritedataReg; // @[mem2wb.scala 107:28]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 88:34]
      RegWriteW <= 1'h0;
    end else if (io_clr) begin // @[mem2wb.scala 88:56]
      RegWriteW <= 1'h0;
    end else if (io_en) begin
      RegWriteW <= io_RegWriteM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 91:34]
      ResultW <= 64'h0;
    end else if (io_clr) begin // @[mem2wb.scala 91:56]
      ResultW <= 64'h0;
    end else if (io_en) begin
      ResultW <= io_ResultM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 92:34]
      WriteRegW <= 5'h0;
    end else if (io_clr) begin // @[mem2wb.scala 92:56]
      WriteRegW <= 5'h0;
    end else if (io_en) begin
      WriteRegW <= io_WriteRegM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 95:34]
      csrWriteW <= 1'h0;
    end else if (io_clr) begin // @[mem2wb.scala 95:56]
      csrWriteW <= 1'h0;
    end else if (io_en) begin
      csrWriteW <= io_csrWriteM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 96:34]
      WritecsrAddrW <= 12'h0;
    end else if (io_clr) begin // @[mem2wb.scala 96:56]
      WritecsrAddrW <= 12'h0;
    end else if (io_en) begin
      WritecsrAddrW <= io_WritecsrAddrM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 98:34]
      PCW <= 64'h0;
    end else if (io_clr) begin // @[mem2wb.scala 98:56]
      PCW <= 64'h0;
    end else if (io_en) begin
      PCW <= io_PCM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 100:34]
      ExceptionTypeW <= 32'h0;
    end else if (io_clr) begin // @[mem2wb.scala 100:56]
      ExceptionTypeW <= 32'h0;
    end else if (io_en) begin
      ExceptionTypeW <= io_ExceptionTypeM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 101:49]
      BranchJump_JrW_Reg <= 2'h0;
    end else if (io_clr) begin // @[mem2wb.scala 101:71]
      BranchJump_JrW_Reg <= 2'h0;
    end else if (io_en) begin
      BranchJump_JrW_Reg <= io_BranchJump_JrM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 103:34]
      ebreak_Reg <= 1'h0;
    end else if (io_clr) begin // @[mem2wb.scala 103:56]
      ebreak_Reg <= 1'h0;
    end else if (io_en) begin
      ebreak_Reg <= io_eBreakM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 104:34]
      pc_nextReg <= 64'h0;
    end else if (io_clr) begin // @[mem2wb.scala 104:56]
      pc_nextReg <= 64'h0;
    end else if (io_en) begin
      pc_nextReg <= io_Pc_NextM;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 105:34]
      Mem_trace_budleReg_pc <= 64'h0;
    end else if (io_clr) begin // @[mem2wb.scala 105:93]
      Mem_trace_budleReg_pc <= 64'h0;
    end else if (io_en) begin
      Mem_trace_budleReg_pc <= io_Mem_trace_budleM_pc;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 105:34]
      Mem_trace_budleReg_data <= 64'h0;
    end else if (io_clr) begin // @[mem2wb.scala 105:93]
      Mem_trace_budleReg_data <= 64'h0;
    end else if (io_en) begin
      Mem_trace_budleReg_data <= io_Mem_trace_budleM_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 105:34]
      Mem_trace_budleReg_mem_fetch_type <= 2'h0;
    end else if (io_clr) begin // @[mem2wb.scala 105:93]
      Mem_trace_budleReg_mem_fetch_type <= 2'h0;
    end else if (io_en) begin
      Mem_trace_budleReg_mem_fetch_type <= io_Mem_trace_budleM_mem_fetch_type;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 105:34]
      Mem_trace_budleReg_addr <= 64'h0;
    end else if (io_clr) begin // @[mem2wb.scala 105:93]
      Mem_trace_budleReg_addr <= 64'h0;
    end else if (io_en) begin
      Mem_trace_budleReg_addr <= io_Mem_trace_budleM_addr;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 105:34]
      Mem_trace_budleReg_len <= 3'h0;
    end else if (io_clr) begin // @[mem2wb.scala 105:93]
      Mem_trace_budleReg_len <= 3'h0;
    end else if (io_en) begin
      Mem_trace_budleReg_len <= io_Mem_trace_budleM_len;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 105:34]
      Mem_trace_budleReg_cache <= 1'h0;
    end else if (io_clr) begin // @[mem2wb.scala 105:93]
      Mem_trace_budleReg_cache <= 1'h0;
    end else if (io_en) begin
      Mem_trace_budleReg_cache <= io_Mem_trace_budleM_cache;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[mem2wb.scala 106:34]
      CsrWritedataReg <= 64'h0;
    end else if (io_clr) begin // @[mem2wb.scala 106:56]
      CsrWritedataReg <= 64'h0;
    end else if (io_en) begin
      CsrWritedataReg <= io_CsrWritedataM;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  RegWriteW = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  ResultW = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  WriteRegW = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  csrWriteW = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  WritecsrAddrW = _RAND_4[11:0];
  _RAND_5 = {2{`RANDOM}};
  PCW = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  ExceptionTypeW = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  BranchJump_JrW_Reg = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  ebreak_Reg = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  pc_nextReg = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  Mem_trace_budleReg_pc = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  Mem_trace_budleReg_data = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  Mem_trace_budleReg_mem_fetch_type = _RAND_12[1:0];
  _RAND_13 = {2{`RANDOM}};
  Mem_trace_budleReg_addr = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  Mem_trace_budleReg_len = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  Mem_trace_budleReg_cache = _RAND_15[0:0];
  _RAND_16 = {2{`RANDOM}};
  CsrWritedataReg = _RAND_16[63:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    RegWriteW = 1'h0;
  end
  if (reset) begin
    ResultW = 64'h0;
  end
  if (reset) begin
    WriteRegW = 5'h0;
  end
  if (reset) begin
    csrWriteW = 1'h0;
  end
  if (reset) begin
    WritecsrAddrW = 12'h0;
  end
  if (reset) begin
    PCW = 64'h0;
  end
  if (reset) begin
    ExceptionTypeW = 32'h0;
  end
  if (reset) begin
    BranchJump_JrW_Reg = 2'h0;
  end
  if (reset) begin
    ebreak_Reg = 1'h0;
  end
  if (reset) begin
    pc_nextReg = 64'h0;
  end
  if (reset) begin
    Mem_trace_budleReg_pc = 64'h0;
  end
  if (reset) begin
    Mem_trace_budleReg_data = 64'h0;
  end
  if (reset) begin
    Mem_trace_budleReg_mem_fetch_type = 2'h0;
  end
  if (reset) begin
    Mem_trace_budleReg_addr = 64'h0;
  end
  if (reset) begin
    Mem_trace_budleReg_len = 3'h0;
  end
  if (reset) begin
    Mem_trace_budleReg_cache = 1'h0;
  end
  if (reset) begin
    CsrWritedataReg = 64'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module addr_cal(
  input  [63:0] io_d_vaddr,
  output [63:0] io_d_paddr,
  output        io_d_cached
);
  assign io_d_paddr = io_d_vaddr; // @[addr_cal.scala 24:16]
  assign io_d_cached = io_d_vaddr[31:29] == 3'h4; // @[macros.scala 479:55]
endmodule
module csa(
  input  [131:0] io_data_0,
  input  [131:0] io_data_1,
  input  [131:0] io_data_2,
  output [131:0] io_result_0,
  output [131:0] io_result_1
);
  wire [131:0] _io_result_0_T = io_data_0 ^ io_data_1; // @[hard_cal.scala 182:32]
  wire [131:0] _io_result_1_T = io_data_0 & io_data_1; // @[hard_cal.scala 183:37]
  wire [131:0] _io_result_1_T_1 = io_data_1 & io_data_2; // @[hard_cal.scala 183:65]
  wire [131:0] _io_result_1_T_2 = _io_result_1_T | _io_result_1_T_1; // @[hard_cal.scala 183:51]
  wire [131:0] _io_result_1_T_3 = io_data_2 & io_data_0; // @[hard_cal.scala 183:93]
  wire [131:0] _io_result_1_T_4 = _io_result_1_T_2 | _io_result_1_T_3; // @[hard_cal.scala 183:79]
  wire [132:0] _io_result_1_T_5 = {_io_result_1_T_4,1'h0}; // @[Cat.scala 31:58]
  assign io_result_0 = _io_result_0_T ^ io_data_2; // @[hard_cal.scala 182:45]
  assign io_result_1 = _io_result_1_T_5[131:0]; // @[hard_cal.scala 183:18]
endmodule
module wallace_adder(
  input          clock,
  input          reset,
  input  [131:0] io_data_in_0,
  input  [131:0] io_data_in_1,
  input  [131:0] io_data_in_2,
  input  [131:0] io_data_in_3,
  input  [131:0] io_data_in_4,
  input  [131:0] io_data_in_5,
  input  [131:0] io_data_in_6,
  input  [131:0] io_data_in_7,
  input  [131:0] io_data_in_8,
  input  [131:0] io_data_in_9,
  input  [131:0] io_data_in_10,
  input  [131:0] io_data_in_11,
  input  [131:0] io_data_in_12,
  input  [131:0] io_data_in_13,
  input  [131:0] io_data_in_14,
  input  [131:0] io_data_in_15,
  input  [131:0] io_data_in_16,
  input  [131:0] io_data_in_17,
  input  [131:0] io_data_in_18,
  input  [131:0] io_data_in_19,
  input  [131:0] io_data_in_20,
  input  [131:0] io_data_in_21,
  input  [131:0] io_data_in_22,
  input  [131:0] io_data_in_23,
  input  [131:0] io_data_in_24,
  input  [131:0] io_data_in_25,
  input  [131:0] io_data_in_26,
  input  [131:0] io_data_in_27,
  input  [131:0] io_data_in_28,
  input  [131:0] io_data_in_29,
  input  [131:0] io_data_in_30,
  input  [131:0] io_data_in_31,
  input  [131:0] io_data_in_32,
  output [131:0] io_result
);
`ifdef RANDOMIZE_REG_INIT
  reg [159:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [159:0] _RAND_4;
  reg [159:0] _RAND_5;
  reg [159:0] _RAND_6;
  reg [159:0] _RAND_7;
  reg [159:0] _RAND_8;
  reg [159:0] _RAND_9;
  reg [159:0] _RAND_10;
  reg [159:0] _RAND_11;
  reg [159:0] _RAND_12;
  reg [159:0] _RAND_13;
  reg [159:0] _RAND_14;
  reg [159:0] _RAND_15;
  reg [159:0] _RAND_16;
  reg [159:0] _RAND_17;
  reg [159:0] _RAND_18;
  reg [159:0] _RAND_19;
  reg [159:0] _RAND_20;
  reg [159:0] _RAND_21;
  reg [159:0] _RAND_22;
  reg [159:0] _RAND_23;
  reg [159:0] _RAND_24;
  reg [159:0] _RAND_25;
  reg [159:0] _RAND_26;
  reg [159:0] _RAND_27;
  reg [159:0] _RAND_28;
  reg [159:0] _RAND_29;
  reg [159:0] _RAND_30;
  reg [159:0] _RAND_31;
  reg [159:0] _RAND_32;
  reg [159:0] _RAND_33;
  reg [159:0] _RAND_34;
  reg [159:0] _RAND_35;
  reg [159:0] _RAND_36;
  reg [159:0] _RAND_37;
  reg [159:0] _RAND_38;
  reg [159:0] _RAND_39;
  reg [159:0] _RAND_40;
  reg [159:0] _RAND_41;
  reg [159:0] _RAND_42;
  reg [159:0] _RAND_43;
  reg [159:0] _RAND_44;
  reg [159:0] _RAND_45;
  reg [159:0] _RAND_46;
  reg [159:0] _RAND_47;
  reg [159:0] _RAND_48;
  reg [159:0] _RAND_49;
  reg [159:0] _RAND_50;
  reg [159:0] _RAND_51;
  reg [159:0] _RAND_52;
  reg [159:0] _RAND_53;
  reg [159:0] _RAND_54;
  reg [159:0] _RAND_55;
  reg [159:0] _RAND_56;
  reg [159:0] _RAND_57;
  reg [159:0] _RAND_58;
  reg [159:0] _RAND_59;
  reg [159:0] _RAND_60;
  reg [159:0] _RAND_61;
  reg [159:0] _RAND_62;
  reg [159:0] _RAND_63;
  reg [159:0] _RAND_64;
  reg [159:0] _RAND_65;
  reg [159:0] _RAND_66;
  reg [159:0] _RAND_67;
`endif // RANDOMIZE_REG_INIT
  wire [131:0] csa_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_1_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_1_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_1_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_1_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_1_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_2_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_2_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_2_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_2_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_2_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_3_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_3_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_3_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_3_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_3_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_4_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_4_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_4_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_4_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_4_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_5_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_5_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_5_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_5_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_5_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_6_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_6_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_6_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_6_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_6_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_7_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_7_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_7_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_7_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_7_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_8_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_8_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_8_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_8_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_8_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_9_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_9_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_9_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_9_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_9_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_10_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_10_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_10_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_10_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_10_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_11_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_11_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_11_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_11_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_11_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_12_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_12_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_12_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_12_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_12_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_13_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_13_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_13_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_13_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_13_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_14_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_14_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_14_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_14_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_14_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_15_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_15_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_15_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_15_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_15_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_16_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_16_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_16_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_16_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_16_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_17_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_17_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_17_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_17_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_17_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_18_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_18_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_18_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_18_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_18_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_19_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_19_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_19_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_19_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_19_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_20_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_20_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_20_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_20_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_20_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_21_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_21_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_21_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_21_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_21_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_22_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_22_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_22_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_22_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_22_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_23_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_23_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_23_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_23_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_23_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_24_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_24_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_24_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_24_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_24_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_25_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_25_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_25_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_25_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_25_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_26_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_26_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_26_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_26_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_26_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_27_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_27_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_27_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_27_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_27_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_28_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_28_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_28_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_28_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_28_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_29_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_29_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_29_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_29_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_29_io_result_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_30_io_data_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_30_io_data_1; // @[hard_cal.scala 204:61]
  wire [131:0] csa_30_io_data_2; // @[hard_cal.scala 204:61]
  wire [131:0] csa_30_io_result_0; // @[hard_cal.scala 204:61]
  wire [131:0] csa_30_io_result_1; // @[hard_cal.scala 204:61]
  reg [131:0] vec_data_out_data_reg__0; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__1; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__2; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__3; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__4; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__5; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__6; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__7; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__8; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__9; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__10; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__11; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__12; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__13; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__14; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__15; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__16; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__17; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__18; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__19; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__20; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg__21; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_1_0; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_1_1; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_1_2; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_1_3; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_1_4; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_1_5; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_1_6; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_1_7; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_1_8; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_1_9; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_1_10; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_1_11; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_1_12; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_1_13; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_1_14; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_2_0; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_2_1; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_2_2; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_2_3; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_2_4; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_2_5; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_2_6; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_2_7; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_2_8; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_2_9; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_3_0; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_3_1; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_3_2; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_3_3; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_3_4; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_3_5; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_3_6; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_4_0; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_4_1; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_4_2; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_4_3; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_4_4; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_5_0; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_5_1; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_5_2; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_5_3; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_6_0; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_6_1; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_out_data_reg_6_2; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_0; // @[hard_cal.scala 220:39]
  reg [131:0] vec_data_1; // @[hard_cal.scala 220:39]
  csa csa ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_io_data_0),
    .io_data_1(csa_io_data_1),
    .io_data_2(csa_io_data_2),
    .io_result_0(csa_io_result_0),
    .io_result_1(csa_io_result_1)
  );
  csa csa_1 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_1_io_data_0),
    .io_data_1(csa_1_io_data_1),
    .io_data_2(csa_1_io_data_2),
    .io_result_0(csa_1_io_result_0),
    .io_result_1(csa_1_io_result_1)
  );
  csa csa_2 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_2_io_data_0),
    .io_data_1(csa_2_io_data_1),
    .io_data_2(csa_2_io_data_2),
    .io_result_0(csa_2_io_result_0),
    .io_result_1(csa_2_io_result_1)
  );
  csa csa_3 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_3_io_data_0),
    .io_data_1(csa_3_io_data_1),
    .io_data_2(csa_3_io_data_2),
    .io_result_0(csa_3_io_result_0),
    .io_result_1(csa_3_io_result_1)
  );
  csa csa_4 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_4_io_data_0),
    .io_data_1(csa_4_io_data_1),
    .io_data_2(csa_4_io_data_2),
    .io_result_0(csa_4_io_result_0),
    .io_result_1(csa_4_io_result_1)
  );
  csa csa_5 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_5_io_data_0),
    .io_data_1(csa_5_io_data_1),
    .io_data_2(csa_5_io_data_2),
    .io_result_0(csa_5_io_result_0),
    .io_result_1(csa_5_io_result_1)
  );
  csa csa_6 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_6_io_data_0),
    .io_data_1(csa_6_io_data_1),
    .io_data_2(csa_6_io_data_2),
    .io_result_0(csa_6_io_result_0),
    .io_result_1(csa_6_io_result_1)
  );
  csa csa_7 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_7_io_data_0),
    .io_data_1(csa_7_io_data_1),
    .io_data_2(csa_7_io_data_2),
    .io_result_0(csa_7_io_result_0),
    .io_result_1(csa_7_io_result_1)
  );
  csa csa_8 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_8_io_data_0),
    .io_data_1(csa_8_io_data_1),
    .io_data_2(csa_8_io_data_2),
    .io_result_0(csa_8_io_result_0),
    .io_result_1(csa_8_io_result_1)
  );
  csa csa_9 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_9_io_data_0),
    .io_data_1(csa_9_io_data_1),
    .io_data_2(csa_9_io_data_2),
    .io_result_0(csa_9_io_result_0),
    .io_result_1(csa_9_io_result_1)
  );
  csa csa_10 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_10_io_data_0),
    .io_data_1(csa_10_io_data_1),
    .io_data_2(csa_10_io_data_2),
    .io_result_0(csa_10_io_result_0),
    .io_result_1(csa_10_io_result_1)
  );
  csa csa_11 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_11_io_data_0),
    .io_data_1(csa_11_io_data_1),
    .io_data_2(csa_11_io_data_2),
    .io_result_0(csa_11_io_result_0),
    .io_result_1(csa_11_io_result_1)
  );
  csa csa_12 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_12_io_data_0),
    .io_data_1(csa_12_io_data_1),
    .io_data_2(csa_12_io_data_2),
    .io_result_0(csa_12_io_result_0),
    .io_result_1(csa_12_io_result_1)
  );
  csa csa_13 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_13_io_data_0),
    .io_data_1(csa_13_io_data_1),
    .io_data_2(csa_13_io_data_2),
    .io_result_0(csa_13_io_result_0),
    .io_result_1(csa_13_io_result_1)
  );
  csa csa_14 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_14_io_data_0),
    .io_data_1(csa_14_io_data_1),
    .io_data_2(csa_14_io_data_2),
    .io_result_0(csa_14_io_result_0),
    .io_result_1(csa_14_io_result_1)
  );
  csa csa_15 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_15_io_data_0),
    .io_data_1(csa_15_io_data_1),
    .io_data_2(csa_15_io_data_2),
    .io_result_0(csa_15_io_result_0),
    .io_result_1(csa_15_io_result_1)
  );
  csa csa_16 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_16_io_data_0),
    .io_data_1(csa_16_io_data_1),
    .io_data_2(csa_16_io_data_2),
    .io_result_0(csa_16_io_result_0),
    .io_result_1(csa_16_io_result_1)
  );
  csa csa_17 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_17_io_data_0),
    .io_data_1(csa_17_io_data_1),
    .io_data_2(csa_17_io_data_2),
    .io_result_0(csa_17_io_result_0),
    .io_result_1(csa_17_io_result_1)
  );
  csa csa_18 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_18_io_data_0),
    .io_data_1(csa_18_io_data_1),
    .io_data_2(csa_18_io_data_2),
    .io_result_0(csa_18_io_result_0),
    .io_result_1(csa_18_io_result_1)
  );
  csa csa_19 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_19_io_data_0),
    .io_data_1(csa_19_io_data_1),
    .io_data_2(csa_19_io_data_2),
    .io_result_0(csa_19_io_result_0),
    .io_result_1(csa_19_io_result_1)
  );
  csa csa_20 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_20_io_data_0),
    .io_data_1(csa_20_io_data_1),
    .io_data_2(csa_20_io_data_2),
    .io_result_0(csa_20_io_result_0),
    .io_result_1(csa_20_io_result_1)
  );
  csa csa_21 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_21_io_data_0),
    .io_data_1(csa_21_io_data_1),
    .io_data_2(csa_21_io_data_2),
    .io_result_0(csa_21_io_result_0),
    .io_result_1(csa_21_io_result_1)
  );
  csa csa_22 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_22_io_data_0),
    .io_data_1(csa_22_io_data_1),
    .io_data_2(csa_22_io_data_2),
    .io_result_0(csa_22_io_result_0),
    .io_result_1(csa_22_io_result_1)
  );
  csa csa_23 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_23_io_data_0),
    .io_data_1(csa_23_io_data_1),
    .io_data_2(csa_23_io_data_2),
    .io_result_0(csa_23_io_result_0),
    .io_result_1(csa_23_io_result_1)
  );
  csa csa_24 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_24_io_data_0),
    .io_data_1(csa_24_io_data_1),
    .io_data_2(csa_24_io_data_2),
    .io_result_0(csa_24_io_result_0),
    .io_result_1(csa_24_io_result_1)
  );
  csa csa_25 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_25_io_data_0),
    .io_data_1(csa_25_io_data_1),
    .io_data_2(csa_25_io_data_2),
    .io_result_0(csa_25_io_result_0),
    .io_result_1(csa_25_io_result_1)
  );
  csa csa_26 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_26_io_data_0),
    .io_data_1(csa_26_io_data_1),
    .io_data_2(csa_26_io_data_2),
    .io_result_0(csa_26_io_result_0),
    .io_result_1(csa_26_io_result_1)
  );
  csa csa_27 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_27_io_data_0),
    .io_data_1(csa_27_io_data_1),
    .io_data_2(csa_27_io_data_2),
    .io_result_0(csa_27_io_result_0),
    .io_result_1(csa_27_io_result_1)
  );
  csa csa_28 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_28_io_data_0),
    .io_data_1(csa_28_io_data_1),
    .io_data_2(csa_28_io_data_2),
    .io_result_0(csa_28_io_result_0),
    .io_result_1(csa_28_io_result_1)
  );
  csa csa_29 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_29_io_data_0),
    .io_data_1(csa_29_io_data_1),
    .io_data_2(csa_29_io_data_2),
    .io_result_0(csa_29_io_result_0),
    .io_result_1(csa_29_io_result_1)
  );
  csa csa_30 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_30_io_data_0),
    .io_data_1(csa_30_io_data_1),
    .io_data_2(csa_30_io_data_2),
    .io_result_0(csa_30_io_result_0),
    .io_result_1(csa_30_io_result_1)
  );
  assign io_result = vec_data_0 + vec_data_1; // @[hard_cal.scala 231:30]
  assign csa_io_data_0 = io_data_in_0; // @[hard_cal.scala 204:36 208:58]
  assign csa_io_data_1 = io_data_in_1; // @[hard_cal.scala 204:36 208:58]
  assign csa_io_data_2 = io_data_in_2; // @[hard_cal.scala 204:36 208:58]
  assign csa_1_io_data_0 = io_data_in_3; // @[hard_cal.scala 204:36 208:58]
  assign csa_1_io_data_1 = io_data_in_4; // @[hard_cal.scala 204:36 208:58]
  assign csa_1_io_data_2 = io_data_in_5; // @[hard_cal.scala 204:36 208:58]
  assign csa_2_io_data_0 = io_data_in_6; // @[hard_cal.scala 204:36 208:58]
  assign csa_2_io_data_1 = io_data_in_7; // @[hard_cal.scala 204:36 208:58]
  assign csa_2_io_data_2 = io_data_in_8; // @[hard_cal.scala 204:36 208:58]
  assign csa_3_io_data_0 = io_data_in_9; // @[hard_cal.scala 204:36 208:58]
  assign csa_3_io_data_1 = io_data_in_10; // @[hard_cal.scala 204:36 208:58]
  assign csa_3_io_data_2 = io_data_in_11; // @[hard_cal.scala 204:36 208:58]
  assign csa_4_io_data_0 = io_data_in_12; // @[hard_cal.scala 204:36 208:58]
  assign csa_4_io_data_1 = io_data_in_13; // @[hard_cal.scala 204:36 208:58]
  assign csa_4_io_data_2 = io_data_in_14; // @[hard_cal.scala 204:36 208:58]
  assign csa_5_io_data_0 = io_data_in_15; // @[hard_cal.scala 204:36 208:58]
  assign csa_5_io_data_1 = io_data_in_16; // @[hard_cal.scala 204:36 208:58]
  assign csa_5_io_data_2 = io_data_in_17; // @[hard_cal.scala 204:36 208:58]
  assign csa_6_io_data_0 = io_data_in_18; // @[hard_cal.scala 204:36 208:58]
  assign csa_6_io_data_1 = io_data_in_19; // @[hard_cal.scala 204:36 208:58]
  assign csa_6_io_data_2 = io_data_in_20; // @[hard_cal.scala 204:36 208:58]
  assign csa_7_io_data_0 = io_data_in_21; // @[hard_cal.scala 204:36 208:58]
  assign csa_7_io_data_1 = io_data_in_22; // @[hard_cal.scala 204:36 208:58]
  assign csa_7_io_data_2 = io_data_in_23; // @[hard_cal.scala 204:36 208:58]
  assign csa_8_io_data_0 = io_data_in_24; // @[hard_cal.scala 204:36 208:58]
  assign csa_8_io_data_1 = io_data_in_25; // @[hard_cal.scala 204:36 208:58]
  assign csa_8_io_data_2 = io_data_in_26; // @[hard_cal.scala 204:36 208:58]
  assign csa_9_io_data_0 = io_data_in_27; // @[hard_cal.scala 204:36 208:58]
  assign csa_9_io_data_1 = io_data_in_28; // @[hard_cal.scala 204:36 208:58]
  assign csa_9_io_data_2 = io_data_in_29; // @[hard_cal.scala 204:36 208:58]
  assign csa_10_io_data_0 = io_data_in_30; // @[hard_cal.scala 204:36 208:58]
  assign csa_10_io_data_1 = io_data_in_31; // @[hard_cal.scala 204:36 208:58]
  assign csa_10_io_data_2 = io_data_in_32; // @[hard_cal.scala 204:36 208:58]
  assign csa_11_io_data_0 = vec_data_out_data_reg__0; // @[hard_cal.scala 204:36 208:58]
  assign csa_11_io_data_1 = vec_data_out_data_reg__1; // @[hard_cal.scala 204:36 208:58]
  assign csa_11_io_data_2 = vec_data_out_data_reg__2; // @[hard_cal.scala 204:36 208:58]
  assign csa_12_io_data_0 = vec_data_out_data_reg__3; // @[hard_cal.scala 204:36 208:58]
  assign csa_12_io_data_1 = vec_data_out_data_reg__4; // @[hard_cal.scala 204:36 208:58]
  assign csa_12_io_data_2 = vec_data_out_data_reg__5; // @[hard_cal.scala 204:36 208:58]
  assign csa_13_io_data_0 = vec_data_out_data_reg__6; // @[hard_cal.scala 204:36 208:58]
  assign csa_13_io_data_1 = vec_data_out_data_reg__7; // @[hard_cal.scala 204:36 208:58]
  assign csa_13_io_data_2 = vec_data_out_data_reg__8; // @[hard_cal.scala 204:36 208:58]
  assign csa_14_io_data_0 = vec_data_out_data_reg__9; // @[hard_cal.scala 204:36 208:58]
  assign csa_14_io_data_1 = vec_data_out_data_reg__10; // @[hard_cal.scala 204:36 208:58]
  assign csa_14_io_data_2 = vec_data_out_data_reg__11; // @[hard_cal.scala 204:36 208:58]
  assign csa_15_io_data_0 = vec_data_out_data_reg__12; // @[hard_cal.scala 204:36 208:58]
  assign csa_15_io_data_1 = vec_data_out_data_reg__13; // @[hard_cal.scala 204:36 208:58]
  assign csa_15_io_data_2 = vec_data_out_data_reg__14; // @[hard_cal.scala 204:36 208:58]
  assign csa_16_io_data_0 = vec_data_out_data_reg__15; // @[hard_cal.scala 204:36 208:58]
  assign csa_16_io_data_1 = vec_data_out_data_reg__16; // @[hard_cal.scala 204:36 208:58]
  assign csa_16_io_data_2 = vec_data_out_data_reg__17; // @[hard_cal.scala 204:36 208:58]
  assign csa_17_io_data_0 = vec_data_out_data_reg__18; // @[hard_cal.scala 204:36 208:58]
  assign csa_17_io_data_1 = vec_data_out_data_reg__19; // @[hard_cal.scala 204:36 208:58]
  assign csa_17_io_data_2 = vec_data_out_data_reg__20; // @[hard_cal.scala 204:36 208:58]
  assign csa_18_io_data_0 = vec_data_out_data_reg_1_0; // @[hard_cal.scala 204:36 208:58]
  assign csa_18_io_data_1 = vec_data_out_data_reg_1_1; // @[hard_cal.scala 204:36 208:58]
  assign csa_18_io_data_2 = vec_data_out_data_reg_1_2; // @[hard_cal.scala 204:36 208:58]
  assign csa_19_io_data_0 = vec_data_out_data_reg_1_3; // @[hard_cal.scala 204:36 208:58]
  assign csa_19_io_data_1 = vec_data_out_data_reg_1_4; // @[hard_cal.scala 204:36 208:58]
  assign csa_19_io_data_2 = vec_data_out_data_reg_1_5; // @[hard_cal.scala 204:36 208:58]
  assign csa_20_io_data_0 = vec_data_out_data_reg_1_6; // @[hard_cal.scala 204:36 208:58]
  assign csa_20_io_data_1 = vec_data_out_data_reg_1_7; // @[hard_cal.scala 204:36 208:58]
  assign csa_20_io_data_2 = vec_data_out_data_reg_1_8; // @[hard_cal.scala 204:36 208:58]
  assign csa_21_io_data_0 = vec_data_out_data_reg_1_9; // @[hard_cal.scala 204:36 208:58]
  assign csa_21_io_data_1 = vec_data_out_data_reg_1_10; // @[hard_cal.scala 204:36 208:58]
  assign csa_21_io_data_2 = vec_data_out_data_reg_1_11; // @[hard_cal.scala 204:36 208:58]
  assign csa_22_io_data_0 = vec_data_out_data_reg_1_12; // @[hard_cal.scala 204:36 208:58]
  assign csa_22_io_data_1 = vec_data_out_data_reg_1_13; // @[hard_cal.scala 204:36 208:58]
  assign csa_22_io_data_2 = vec_data_out_data_reg_1_14; // @[hard_cal.scala 204:36 208:58]
  assign csa_23_io_data_0 = vec_data_out_data_reg_2_0; // @[hard_cal.scala 204:36 208:58]
  assign csa_23_io_data_1 = vec_data_out_data_reg_2_1; // @[hard_cal.scala 204:36 208:58]
  assign csa_23_io_data_2 = vec_data_out_data_reg_2_2; // @[hard_cal.scala 204:36 208:58]
  assign csa_24_io_data_0 = vec_data_out_data_reg_2_3; // @[hard_cal.scala 204:36 208:58]
  assign csa_24_io_data_1 = vec_data_out_data_reg_2_4; // @[hard_cal.scala 204:36 208:58]
  assign csa_24_io_data_2 = vec_data_out_data_reg_2_5; // @[hard_cal.scala 204:36 208:58]
  assign csa_25_io_data_0 = vec_data_out_data_reg_2_6; // @[hard_cal.scala 204:36 208:58]
  assign csa_25_io_data_1 = vec_data_out_data_reg_2_7; // @[hard_cal.scala 204:36 208:58]
  assign csa_25_io_data_2 = vec_data_out_data_reg_2_8; // @[hard_cal.scala 204:36 208:58]
  assign csa_26_io_data_0 = vec_data_out_data_reg_3_0; // @[hard_cal.scala 204:36 208:58]
  assign csa_26_io_data_1 = vec_data_out_data_reg_3_1; // @[hard_cal.scala 204:36 208:58]
  assign csa_26_io_data_2 = vec_data_out_data_reg_3_2; // @[hard_cal.scala 204:36 208:58]
  assign csa_27_io_data_0 = vec_data_out_data_reg_3_3; // @[hard_cal.scala 204:36 208:58]
  assign csa_27_io_data_1 = vec_data_out_data_reg_3_4; // @[hard_cal.scala 204:36 208:58]
  assign csa_27_io_data_2 = vec_data_out_data_reg_3_5; // @[hard_cal.scala 204:36 208:58]
  assign csa_28_io_data_0 = vec_data_out_data_reg_4_0; // @[hard_cal.scala 204:36 208:58]
  assign csa_28_io_data_1 = vec_data_out_data_reg_4_1; // @[hard_cal.scala 204:36 208:58]
  assign csa_28_io_data_2 = vec_data_out_data_reg_4_2; // @[hard_cal.scala 204:36 208:58]
  assign csa_29_io_data_0 = vec_data_out_data_reg_5_0; // @[hard_cal.scala 204:36 208:58]
  assign csa_29_io_data_1 = vec_data_out_data_reg_5_1; // @[hard_cal.scala 204:36 208:58]
  assign csa_29_io_data_2 = vec_data_out_data_reg_5_2; // @[hard_cal.scala 204:36 208:58]
  assign csa_30_io_data_0 = vec_data_out_data_reg_6_0; // @[hard_cal.scala 204:36 208:58]
  assign csa_30_io_data_1 = vec_data_out_data_reg_6_1; // @[hard_cal.scala 204:36 208:58]
  assign csa_30_io_data_2 = vec_data_out_data_reg_6_2; // @[hard_cal.scala 204:36 208:58]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__0 <= 132'h0;
    end else begin
      vec_data_out_data_reg__0 <= csa_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__1 <= 132'h0;
    end else begin
      vec_data_out_data_reg__1 <= csa_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__2 <= 132'h0;
    end else begin
      vec_data_out_data_reg__2 <= csa_1_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__3 <= 132'h0;
    end else begin
      vec_data_out_data_reg__3 <= csa_1_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__4 <= 132'h0;
    end else begin
      vec_data_out_data_reg__4 <= csa_2_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__5 <= 132'h0;
    end else begin
      vec_data_out_data_reg__5 <= csa_2_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__6 <= 132'h0;
    end else begin
      vec_data_out_data_reg__6 <= csa_3_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__7 <= 132'h0;
    end else begin
      vec_data_out_data_reg__7 <= csa_3_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__8 <= 132'h0;
    end else begin
      vec_data_out_data_reg__8 <= csa_4_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__9 <= 132'h0;
    end else begin
      vec_data_out_data_reg__9 <= csa_4_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__10 <= 132'h0;
    end else begin
      vec_data_out_data_reg__10 <= csa_5_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__11 <= 132'h0;
    end else begin
      vec_data_out_data_reg__11 <= csa_5_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__12 <= 132'h0;
    end else begin
      vec_data_out_data_reg__12 <= csa_6_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__13 <= 132'h0;
    end else begin
      vec_data_out_data_reg__13 <= csa_6_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__14 <= 132'h0;
    end else begin
      vec_data_out_data_reg__14 <= csa_7_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__15 <= 132'h0;
    end else begin
      vec_data_out_data_reg__15 <= csa_7_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__16 <= 132'h0;
    end else begin
      vec_data_out_data_reg__16 <= csa_8_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__17 <= 132'h0;
    end else begin
      vec_data_out_data_reg__17 <= csa_8_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__18 <= 132'h0;
    end else begin
      vec_data_out_data_reg__18 <= csa_9_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__19 <= 132'h0;
    end else begin
      vec_data_out_data_reg__19 <= csa_9_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__20 <= 132'h0;
    end else begin
      vec_data_out_data_reg__20 <= csa_10_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__21 <= 132'h0;
    end else begin
      vec_data_out_data_reg__21 <= csa_10_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_0 <= 132'h0;
    end else begin
      vec_data_out_data_reg_1_0 <= csa_11_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_1 <= 132'h0;
    end else begin
      vec_data_out_data_reg_1_1 <= csa_11_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_2 <= 132'h0;
    end else begin
      vec_data_out_data_reg_1_2 <= csa_12_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_3 <= 132'h0;
    end else begin
      vec_data_out_data_reg_1_3 <= csa_12_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_4 <= 132'h0;
    end else begin
      vec_data_out_data_reg_1_4 <= csa_13_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_5 <= 132'h0;
    end else begin
      vec_data_out_data_reg_1_5 <= csa_13_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_6 <= 132'h0;
    end else begin
      vec_data_out_data_reg_1_6 <= csa_14_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_7 <= 132'h0;
    end else begin
      vec_data_out_data_reg_1_7 <= csa_14_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_8 <= 132'h0;
    end else begin
      vec_data_out_data_reg_1_8 <= csa_15_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_9 <= 132'h0;
    end else begin
      vec_data_out_data_reg_1_9 <= csa_15_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_10 <= 132'h0;
    end else begin
      vec_data_out_data_reg_1_10 <= csa_16_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_11 <= 132'h0;
    end else begin
      vec_data_out_data_reg_1_11 <= csa_16_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_12 <= 132'h0;
    end else begin
      vec_data_out_data_reg_1_12 <= csa_17_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_13 <= 132'h0;
    end else begin
      vec_data_out_data_reg_1_13 <= csa_17_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 211:39 217:44]
      vec_data_out_data_reg_1_14 <= 132'h0;
    end else begin
      vec_data_out_data_reg_1_14 <= vec_data_out_data_reg__21;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_2_0 <= 132'h0;
    end else begin
      vec_data_out_data_reg_2_0 <= csa_18_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_2_1 <= 132'h0;
    end else begin
      vec_data_out_data_reg_2_1 <= csa_18_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_2_2 <= 132'h0;
    end else begin
      vec_data_out_data_reg_2_2 <= csa_19_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_2_3 <= 132'h0;
    end else begin
      vec_data_out_data_reg_2_3 <= csa_19_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_2_4 <= 132'h0;
    end else begin
      vec_data_out_data_reg_2_4 <= csa_20_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_2_5 <= 132'h0;
    end else begin
      vec_data_out_data_reg_2_5 <= csa_20_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_2_6 <= 132'h0;
    end else begin
      vec_data_out_data_reg_2_6 <= csa_21_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_2_7 <= 132'h0;
    end else begin
      vec_data_out_data_reg_2_7 <= csa_21_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_2_8 <= 132'h0;
    end else begin
      vec_data_out_data_reg_2_8 <= csa_22_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_2_9 <= 132'h0;
    end else begin
      vec_data_out_data_reg_2_9 <= csa_22_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_3_0 <= 132'h0;
    end else begin
      vec_data_out_data_reg_3_0 <= csa_23_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_3_1 <= 132'h0;
    end else begin
      vec_data_out_data_reg_3_1 <= csa_23_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_3_2 <= 132'h0;
    end else begin
      vec_data_out_data_reg_3_2 <= csa_24_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_3_3 <= 132'h0;
    end else begin
      vec_data_out_data_reg_3_3 <= csa_24_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_3_4 <= 132'h0;
    end else begin
      vec_data_out_data_reg_3_4 <= csa_25_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_3_5 <= 132'h0;
    end else begin
      vec_data_out_data_reg_3_5 <= csa_25_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 211:39 217:44]
      vec_data_out_data_reg_3_6 <= 132'h0;
    end else begin
      vec_data_out_data_reg_3_6 <= vec_data_out_data_reg_2_9;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_4_0 <= 132'h0;
    end else begin
      vec_data_out_data_reg_4_0 <= csa_26_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_4_1 <= 132'h0;
    end else begin
      vec_data_out_data_reg_4_1 <= csa_26_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_4_2 <= 132'h0;
    end else begin
      vec_data_out_data_reg_4_2 <= csa_27_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_4_3 <= 132'h0;
    end else begin
      vec_data_out_data_reg_4_3 <= csa_27_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 211:39 217:44]
      vec_data_out_data_reg_4_4 <= 132'h0;
    end else begin
      vec_data_out_data_reg_4_4 <= vec_data_out_data_reg_3_6;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_5_0 <= 132'h0;
    end else begin
      vec_data_out_data_reg_5_0 <= csa_28_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_5_1 <= 132'h0;
    end else begin
      vec_data_out_data_reg_5_1 <= csa_28_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 211:39 217:44]
      vec_data_out_data_reg_5_2 <= 132'h0;
    end else begin
      vec_data_out_data_reg_5_2 <= vec_data_out_data_reg_4_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 211:39 217:44]
      vec_data_out_data_reg_5_3 <= 132'h0;
    end else begin
      vec_data_out_data_reg_5_3 <= vec_data_out_data_reg_4_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_6_0 <= 132'h0;
    end else begin
      vec_data_out_data_reg_6_0 <= csa_29_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_6_1 <= 132'h0;
    end else begin
      vec_data_out_data_reg_6_1 <= csa_29_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 211:39 217:44]
      vec_data_out_data_reg_6_2 <= 132'h0;
    end else begin
      vec_data_out_data_reg_6_2 <= vec_data_out_data_reg_5_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_0 <= 132'h0;
    end else begin
      vec_data_0 <= csa_30_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_1 <= 132'h0;
    end else begin
      vec_data_1 <= csa_30_io_result_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {5{`RANDOM}};
  vec_data_out_data_reg__0 = _RAND_0[131:0];
  _RAND_1 = {5{`RANDOM}};
  vec_data_out_data_reg__1 = _RAND_1[131:0];
  _RAND_2 = {5{`RANDOM}};
  vec_data_out_data_reg__2 = _RAND_2[131:0];
  _RAND_3 = {5{`RANDOM}};
  vec_data_out_data_reg__3 = _RAND_3[131:0];
  _RAND_4 = {5{`RANDOM}};
  vec_data_out_data_reg__4 = _RAND_4[131:0];
  _RAND_5 = {5{`RANDOM}};
  vec_data_out_data_reg__5 = _RAND_5[131:0];
  _RAND_6 = {5{`RANDOM}};
  vec_data_out_data_reg__6 = _RAND_6[131:0];
  _RAND_7 = {5{`RANDOM}};
  vec_data_out_data_reg__7 = _RAND_7[131:0];
  _RAND_8 = {5{`RANDOM}};
  vec_data_out_data_reg__8 = _RAND_8[131:0];
  _RAND_9 = {5{`RANDOM}};
  vec_data_out_data_reg__9 = _RAND_9[131:0];
  _RAND_10 = {5{`RANDOM}};
  vec_data_out_data_reg__10 = _RAND_10[131:0];
  _RAND_11 = {5{`RANDOM}};
  vec_data_out_data_reg__11 = _RAND_11[131:0];
  _RAND_12 = {5{`RANDOM}};
  vec_data_out_data_reg__12 = _RAND_12[131:0];
  _RAND_13 = {5{`RANDOM}};
  vec_data_out_data_reg__13 = _RAND_13[131:0];
  _RAND_14 = {5{`RANDOM}};
  vec_data_out_data_reg__14 = _RAND_14[131:0];
  _RAND_15 = {5{`RANDOM}};
  vec_data_out_data_reg__15 = _RAND_15[131:0];
  _RAND_16 = {5{`RANDOM}};
  vec_data_out_data_reg__16 = _RAND_16[131:0];
  _RAND_17 = {5{`RANDOM}};
  vec_data_out_data_reg__17 = _RAND_17[131:0];
  _RAND_18 = {5{`RANDOM}};
  vec_data_out_data_reg__18 = _RAND_18[131:0];
  _RAND_19 = {5{`RANDOM}};
  vec_data_out_data_reg__19 = _RAND_19[131:0];
  _RAND_20 = {5{`RANDOM}};
  vec_data_out_data_reg__20 = _RAND_20[131:0];
  _RAND_21 = {5{`RANDOM}};
  vec_data_out_data_reg__21 = _RAND_21[131:0];
  _RAND_22 = {5{`RANDOM}};
  vec_data_out_data_reg_1_0 = _RAND_22[131:0];
  _RAND_23 = {5{`RANDOM}};
  vec_data_out_data_reg_1_1 = _RAND_23[131:0];
  _RAND_24 = {5{`RANDOM}};
  vec_data_out_data_reg_1_2 = _RAND_24[131:0];
  _RAND_25 = {5{`RANDOM}};
  vec_data_out_data_reg_1_3 = _RAND_25[131:0];
  _RAND_26 = {5{`RANDOM}};
  vec_data_out_data_reg_1_4 = _RAND_26[131:0];
  _RAND_27 = {5{`RANDOM}};
  vec_data_out_data_reg_1_5 = _RAND_27[131:0];
  _RAND_28 = {5{`RANDOM}};
  vec_data_out_data_reg_1_6 = _RAND_28[131:0];
  _RAND_29 = {5{`RANDOM}};
  vec_data_out_data_reg_1_7 = _RAND_29[131:0];
  _RAND_30 = {5{`RANDOM}};
  vec_data_out_data_reg_1_8 = _RAND_30[131:0];
  _RAND_31 = {5{`RANDOM}};
  vec_data_out_data_reg_1_9 = _RAND_31[131:0];
  _RAND_32 = {5{`RANDOM}};
  vec_data_out_data_reg_1_10 = _RAND_32[131:0];
  _RAND_33 = {5{`RANDOM}};
  vec_data_out_data_reg_1_11 = _RAND_33[131:0];
  _RAND_34 = {5{`RANDOM}};
  vec_data_out_data_reg_1_12 = _RAND_34[131:0];
  _RAND_35 = {5{`RANDOM}};
  vec_data_out_data_reg_1_13 = _RAND_35[131:0];
  _RAND_36 = {5{`RANDOM}};
  vec_data_out_data_reg_1_14 = _RAND_36[131:0];
  _RAND_37 = {5{`RANDOM}};
  vec_data_out_data_reg_2_0 = _RAND_37[131:0];
  _RAND_38 = {5{`RANDOM}};
  vec_data_out_data_reg_2_1 = _RAND_38[131:0];
  _RAND_39 = {5{`RANDOM}};
  vec_data_out_data_reg_2_2 = _RAND_39[131:0];
  _RAND_40 = {5{`RANDOM}};
  vec_data_out_data_reg_2_3 = _RAND_40[131:0];
  _RAND_41 = {5{`RANDOM}};
  vec_data_out_data_reg_2_4 = _RAND_41[131:0];
  _RAND_42 = {5{`RANDOM}};
  vec_data_out_data_reg_2_5 = _RAND_42[131:0];
  _RAND_43 = {5{`RANDOM}};
  vec_data_out_data_reg_2_6 = _RAND_43[131:0];
  _RAND_44 = {5{`RANDOM}};
  vec_data_out_data_reg_2_7 = _RAND_44[131:0];
  _RAND_45 = {5{`RANDOM}};
  vec_data_out_data_reg_2_8 = _RAND_45[131:0];
  _RAND_46 = {5{`RANDOM}};
  vec_data_out_data_reg_2_9 = _RAND_46[131:0];
  _RAND_47 = {5{`RANDOM}};
  vec_data_out_data_reg_3_0 = _RAND_47[131:0];
  _RAND_48 = {5{`RANDOM}};
  vec_data_out_data_reg_3_1 = _RAND_48[131:0];
  _RAND_49 = {5{`RANDOM}};
  vec_data_out_data_reg_3_2 = _RAND_49[131:0];
  _RAND_50 = {5{`RANDOM}};
  vec_data_out_data_reg_3_3 = _RAND_50[131:0];
  _RAND_51 = {5{`RANDOM}};
  vec_data_out_data_reg_3_4 = _RAND_51[131:0];
  _RAND_52 = {5{`RANDOM}};
  vec_data_out_data_reg_3_5 = _RAND_52[131:0];
  _RAND_53 = {5{`RANDOM}};
  vec_data_out_data_reg_3_6 = _RAND_53[131:0];
  _RAND_54 = {5{`RANDOM}};
  vec_data_out_data_reg_4_0 = _RAND_54[131:0];
  _RAND_55 = {5{`RANDOM}};
  vec_data_out_data_reg_4_1 = _RAND_55[131:0];
  _RAND_56 = {5{`RANDOM}};
  vec_data_out_data_reg_4_2 = _RAND_56[131:0];
  _RAND_57 = {5{`RANDOM}};
  vec_data_out_data_reg_4_3 = _RAND_57[131:0];
  _RAND_58 = {5{`RANDOM}};
  vec_data_out_data_reg_4_4 = _RAND_58[131:0];
  _RAND_59 = {5{`RANDOM}};
  vec_data_out_data_reg_5_0 = _RAND_59[131:0];
  _RAND_60 = {5{`RANDOM}};
  vec_data_out_data_reg_5_1 = _RAND_60[131:0];
  _RAND_61 = {5{`RANDOM}};
  vec_data_out_data_reg_5_2 = _RAND_61[131:0];
  _RAND_62 = {5{`RANDOM}};
  vec_data_out_data_reg_5_3 = _RAND_62[131:0];
  _RAND_63 = {5{`RANDOM}};
  vec_data_out_data_reg_6_0 = _RAND_63[131:0];
  _RAND_64 = {5{`RANDOM}};
  vec_data_out_data_reg_6_1 = _RAND_64[131:0];
  _RAND_65 = {5{`RANDOM}};
  vec_data_out_data_reg_6_2 = _RAND_65[131:0];
  _RAND_66 = {5{`RANDOM}};
  vec_data_0 = _RAND_66[131:0];
  _RAND_67 = {5{`RANDOM}};
  vec_data_1 = _RAND_67[131:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    vec_data_out_data_reg__0 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__1 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__2 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__3 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__4 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__5 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__6 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__7 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__8 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__9 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__10 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__11 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__12 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__13 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__14 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__15 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__16 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__17 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__18 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__19 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__20 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__21 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_0 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_1 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_2 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_3 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_4 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_5 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_6 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_7 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_8 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_9 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_10 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_11 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_12 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_13 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_14 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_2_0 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_2_1 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_2_2 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_2_3 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_2_4 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_2_5 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_2_6 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_2_7 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_2_8 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_2_9 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_3_0 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_3_1 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_3_2 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_3_3 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_3_4 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_3_5 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_3_6 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_4_0 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_4_1 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_4_2 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_4_3 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_4_4 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_5_0 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_5_1 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_5_2 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_5_3 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_6_0 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_6_1 = 132'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_6_2 = 132'h0;
  end
  if (reset) begin
    vec_data_0 = 132'h0;
  end
  if (reset) begin
    vec_data_1 = 132'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module mul_hard(
  input         clock,
  input         reset,
  output [65:0] io_result_0,
  output [65:0] io_result_1,
  input  [65:0] io_data_0,
  input  [65:0] io_data_1,
  input         io_input_valid,
  output        io_input_ready,
  output        io_Output_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [159:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [159:0] _RAND_4;
  reg [159:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  cal_module_clock; // @[hard_cal.scala 295:28]
  wire  cal_module_reset; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_0; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_1; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_2; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_3; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_4; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_5; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_6; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_7; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_8; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_9; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_10; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_11; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_12; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_13; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_14; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_15; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_16; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_17; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_18; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_19; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_20; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_21; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_22; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_23; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_24; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_25; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_26; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_27; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_28; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_29; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_30; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_31; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_data_in_32; // @[hard_cal.scala 295:28]
  wire [131:0] cal_module_io_result; // @[hard_cal.scala 295:28]
  reg [131:0] regs_0; // @[hard_cal.scala 254:23]
  reg [131:0] regs_1; // @[hard_cal.scala 254:23]
  reg [6:0] counter; // @[hard_cal.scala 256:26]
  reg  cal_start; // @[hard_cal.scala 257:28]
  wire [6:0] _counter_T_1 = counter + 7'h1; // @[hard_cal.scala 259:39]
  wire  _signed_T = io_input_valid & io_input_ready; // @[hard_cal.scala 260:35]
  reg [131:0] result_reg; // @[hard_cal.scala 261:29]
  reg [131:0] x_fu; // @[hard_cal.scala 264:23]
  wire [2:0] look_up_data = {regs_1[1],regs_1[0],1'h0}; // @[Cat.scala 31:58]
  wire [132:0] _booth_data_0_T = {regs_0, 1'h0}; // @[hard_cal.scala 279:38]
  wire [132:0] _booth_data_0_T_1 = {x_fu, 1'h0}; // @[hard_cal.scala 280:31]
  wire [131:0] _booth_data_0_T_3 = 3'h1 == look_up_data ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_0_T_5 = 3'h2 == look_up_data ? regs_0 : _booth_data_0_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_0_T_7 = 3'h3 == look_up_data ? _booth_data_0_T : {{1'd0}, _booth_data_0_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_0_T_9 = 3'h4 == look_up_data ? _booth_data_0_T_1 : _booth_data_0_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_0_T_11 = 3'h5 == look_up_data ? {{1'd0}, x_fu} : _booth_data_0_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_0_T_13 = 3'h6 == look_up_data ? {{1'd0}, x_fu} : _booth_data_0_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_0_T_15 = 3'h7 == look_up_data ? 133'h0 : _booth_data_0_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_0_T_17 = {1'h0,_booth_data_0_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_0_T_18 = {{1'd0}, _booth_data_0_T_17}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_1 = {regs_1[3],regs_1[2],regs_1[1]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_1_T_3 = 3'h1 == look_up_data_1 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_1_T_5 = 3'h2 == look_up_data_1 ? regs_0 : _booth_data_1_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_1_T_7 = 3'h3 == look_up_data_1 ? _booth_data_0_T : {{1'd0}, _booth_data_1_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_1_T_9 = 3'h4 == look_up_data_1 ? _booth_data_0_T_1 : _booth_data_1_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_1_T_11 = 3'h5 == look_up_data_1 ? {{1'd0}, x_fu} : _booth_data_1_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_1_T_13 = 3'h6 == look_up_data_1 ? {{1'd0}, x_fu} : _booth_data_1_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_1_T_15 = 3'h7 == look_up_data_1 ? 133'h0 : _booth_data_1_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_1_T_17 = {1'h0,_booth_data_1_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [68:0] _GEN_0 = {_booth_data_1_T_17, 2'h0}; // @[hard_cal.scala 285:19]
  wire [69:0] _booth_data_1_T_18 = {{1'd0}, _GEN_0}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_2 = {regs_1[5],regs_1[4],regs_1[3]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_2_T_3 = 3'h1 == look_up_data_2 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_2_T_5 = 3'h2 == look_up_data_2 ? regs_0 : _booth_data_2_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_2_T_7 = 3'h3 == look_up_data_2 ? _booth_data_0_T : {{1'd0}, _booth_data_2_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_2_T_9 = 3'h4 == look_up_data_2 ? _booth_data_0_T_1 : _booth_data_2_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_2_T_11 = 3'h5 == look_up_data_2 ? {{1'd0}, x_fu} : _booth_data_2_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_2_T_13 = 3'h6 == look_up_data_2 ? {{1'd0}, x_fu} : _booth_data_2_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_2_T_15 = 3'h7 == look_up_data_2 ? 133'h0 : _booth_data_2_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_2_T_17 = {1'h0,_booth_data_2_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [70:0] _GEN_1 = {_booth_data_2_T_17, 4'h0}; // @[hard_cal.scala 285:19]
  wire [73:0] _booth_data_2_T_18 = {{3'd0}, _GEN_1}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_3 = {regs_1[7],regs_1[6],regs_1[5]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_3_T_3 = 3'h1 == look_up_data_3 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_3_T_5 = 3'h2 == look_up_data_3 ? regs_0 : _booth_data_3_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_3_T_7 = 3'h3 == look_up_data_3 ? _booth_data_0_T : {{1'd0}, _booth_data_3_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_3_T_9 = 3'h4 == look_up_data_3 ? _booth_data_0_T_1 : _booth_data_3_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_3_T_11 = 3'h5 == look_up_data_3 ? {{1'd0}, x_fu} : _booth_data_3_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_3_T_13 = 3'h6 == look_up_data_3 ? {{1'd0}, x_fu} : _booth_data_3_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_3_T_15 = 3'h7 == look_up_data_3 ? 133'h0 : _booth_data_3_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_3_T_17 = {1'h0,_booth_data_3_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [72:0] _GEN_2 = {_booth_data_3_T_17, 6'h0}; // @[hard_cal.scala 285:19]
  wire [73:0] _booth_data_3_T_18 = {{1'd0}, _GEN_2}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_4 = {regs_1[9],regs_1[8],regs_1[7]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_4_T_3 = 3'h1 == look_up_data_4 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_4_T_5 = 3'h2 == look_up_data_4 ? regs_0 : _booth_data_4_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_4_T_7 = 3'h3 == look_up_data_4 ? _booth_data_0_T : {{1'd0}, _booth_data_4_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_4_T_9 = 3'h4 == look_up_data_4 ? _booth_data_0_T_1 : _booth_data_4_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_4_T_11 = 3'h5 == look_up_data_4 ? {{1'd0}, x_fu} : _booth_data_4_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_4_T_13 = 3'h6 == look_up_data_4 ? {{1'd0}, x_fu} : _booth_data_4_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_4_T_15 = 3'h7 == look_up_data_4 ? 133'h0 : _booth_data_4_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_4_T_17 = {1'h0,_booth_data_4_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [74:0] _GEN_3 = {_booth_data_4_T_17, 8'h0}; // @[hard_cal.scala 285:19]
  wire [81:0] _booth_data_4_T_18 = {{7'd0}, _GEN_3}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_5 = {regs_1[11],regs_1[10],regs_1[9]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_5_T_3 = 3'h1 == look_up_data_5 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_5_T_5 = 3'h2 == look_up_data_5 ? regs_0 : _booth_data_5_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_5_T_7 = 3'h3 == look_up_data_5 ? _booth_data_0_T : {{1'd0}, _booth_data_5_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_5_T_9 = 3'h4 == look_up_data_5 ? _booth_data_0_T_1 : _booth_data_5_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_5_T_11 = 3'h5 == look_up_data_5 ? {{1'd0}, x_fu} : _booth_data_5_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_5_T_13 = 3'h6 == look_up_data_5 ? {{1'd0}, x_fu} : _booth_data_5_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_5_T_15 = 3'h7 == look_up_data_5 ? 133'h0 : _booth_data_5_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_5_T_17 = {1'h0,_booth_data_5_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [76:0] _GEN_4 = {_booth_data_5_T_17, 10'h0}; // @[hard_cal.scala 285:19]
  wire [81:0] _booth_data_5_T_18 = {{5'd0}, _GEN_4}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_6 = {regs_1[13],regs_1[12],regs_1[11]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_6_T_3 = 3'h1 == look_up_data_6 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_6_T_5 = 3'h2 == look_up_data_6 ? regs_0 : _booth_data_6_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_6_T_7 = 3'h3 == look_up_data_6 ? _booth_data_0_T : {{1'd0}, _booth_data_6_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_6_T_9 = 3'h4 == look_up_data_6 ? _booth_data_0_T_1 : _booth_data_6_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_6_T_11 = 3'h5 == look_up_data_6 ? {{1'd0}, x_fu} : _booth_data_6_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_6_T_13 = 3'h6 == look_up_data_6 ? {{1'd0}, x_fu} : _booth_data_6_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_6_T_15 = 3'h7 == look_up_data_6 ? 133'h0 : _booth_data_6_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_6_T_17 = {1'h0,_booth_data_6_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [78:0] _GEN_5 = {_booth_data_6_T_17, 12'h0}; // @[hard_cal.scala 285:19]
  wire [81:0] _booth_data_6_T_18 = {{3'd0}, _GEN_5}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_7 = {regs_1[15],regs_1[14],regs_1[13]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_7_T_3 = 3'h1 == look_up_data_7 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_7_T_5 = 3'h2 == look_up_data_7 ? regs_0 : _booth_data_7_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_7_T_7 = 3'h3 == look_up_data_7 ? _booth_data_0_T : {{1'd0}, _booth_data_7_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_7_T_9 = 3'h4 == look_up_data_7 ? _booth_data_0_T_1 : _booth_data_7_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_7_T_11 = 3'h5 == look_up_data_7 ? {{1'd0}, x_fu} : _booth_data_7_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_7_T_13 = 3'h6 == look_up_data_7 ? {{1'd0}, x_fu} : _booth_data_7_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_7_T_15 = 3'h7 == look_up_data_7 ? 133'h0 : _booth_data_7_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_7_T_17 = {1'h0,_booth_data_7_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [80:0] _GEN_6 = {_booth_data_7_T_17, 14'h0}; // @[hard_cal.scala 285:19]
  wire [81:0] _booth_data_7_T_18 = {{1'd0}, _GEN_6}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_8 = {regs_1[17],regs_1[16],regs_1[15]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_8_T_3 = 3'h1 == look_up_data_8 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_8_T_5 = 3'h2 == look_up_data_8 ? regs_0 : _booth_data_8_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_8_T_7 = 3'h3 == look_up_data_8 ? _booth_data_0_T : {{1'd0}, _booth_data_8_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_8_T_9 = 3'h4 == look_up_data_8 ? _booth_data_0_T_1 : _booth_data_8_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_8_T_11 = 3'h5 == look_up_data_8 ? {{1'd0}, x_fu} : _booth_data_8_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_8_T_13 = 3'h6 == look_up_data_8 ? {{1'd0}, x_fu} : _booth_data_8_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_8_T_15 = 3'h7 == look_up_data_8 ? 133'h0 : _booth_data_8_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_8_T_17 = {1'h0,_booth_data_8_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [82:0] _GEN_7 = {_booth_data_8_T_17, 16'h0}; // @[hard_cal.scala 285:19]
  wire [97:0] _booth_data_8_T_18 = {{15'd0}, _GEN_7}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_9 = {regs_1[19],regs_1[18],regs_1[17]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_9_T_3 = 3'h1 == look_up_data_9 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_9_T_5 = 3'h2 == look_up_data_9 ? regs_0 : _booth_data_9_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_9_T_7 = 3'h3 == look_up_data_9 ? _booth_data_0_T : {{1'd0}, _booth_data_9_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_9_T_9 = 3'h4 == look_up_data_9 ? _booth_data_0_T_1 : _booth_data_9_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_9_T_11 = 3'h5 == look_up_data_9 ? {{1'd0}, x_fu} : _booth_data_9_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_9_T_13 = 3'h6 == look_up_data_9 ? {{1'd0}, x_fu} : _booth_data_9_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_9_T_15 = 3'h7 == look_up_data_9 ? 133'h0 : _booth_data_9_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_9_T_17 = {1'h0,_booth_data_9_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [84:0] _GEN_8 = {_booth_data_9_T_17, 18'h0}; // @[hard_cal.scala 285:19]
  wire [97:0] _booth_data_9_T_18 = {{13'd0}, _GEN_8}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_10 = {regs_1[21],regs_1[20],regs_1[19]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_10_T_3 = 3'h1 == look_up_data_10 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_10_T_5 = 3'h2 == look_up_data_10 ? regs_0 : _booth_data_10_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_10_T_7 = 3'h3 == look_up_data_10 ? _booth_data_0_T : {{1'd0}, _booth_data_10_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_10_T_9 = 3'h4 == look_up_data_10 ? _booth_data_0_T_1 : _booth_data_10_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_10_T_11 = 3'h5 == look_up_data_10 ? {{1'd0}, x_fu} : _booth_data_10_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_10_T_13 = 3'h6 == look_up_data_10 ? {{1'd0}, x_fu} : _booth_data_10_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_10_T_15 = 3'h7 == look_up_data_10 ? 133'h0 : _booth_data_10_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_10_T_17 = {1'h0,_booth_data_10_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [86:0] _GEN_9 = {_booth_data_10_T_17, 20'h0}; // @[hard_cal.scala 285:19]
  wire [97:0] _booth_data_10_T_18 = {{11'd0}, _GEN_9}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_11 = {regs_1[23],regs_1[22],regs_1[21]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_11_T_3 = 3'h1 == look_up_data_11 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_11_T_5 = 3'h2 == look_up_data_11 ? regs_0 : _booth_data_11_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_11_T_7 = 3'h3 == look_up_data_11 ? _booth_data_0_T : {{1'd0}, _booth_data_11_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_11_T_9 = 3'h4 == look_up_data_11 ? _booth_data_0_T_1 : _booth_data_11_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_11_T_11 = 3'h5 == look_up_data_11 ? {{1'd0}, x_fu} : _booth_data_11_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_11_T_13 = 3'h6 == look_up_data_11 ? {{1'd0}, x_fu} : _booth_data_11_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_11_T_15 = 3'h7 == look_up_data_11 ? 133'h0 : _booth_data_11_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_11_T_17 = {1'h0,_booth_data_11_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [88:0] _GEN_10 = {_booth_data_11_T_17, 22'h0}; // @[hard_cal.scala 285:19]
  wire [97:0] _booth_data_11_T_18 = {{9'd0}, _GEN_10}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_12 = {regs_1[25],regs_1[24],regs_1[23]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_12_T_3 = 3'h1 == look_up_data_12 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_12_T_5 = 3'h2 == look_up_data_12 ? regs_0 : _booth_data_12_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_12_T_7 = 3'h3 == look_up_data_12 ? _booth_data_0_T : {{1'd0}, _booth_data_12_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_12_T_9 = 3'h4 == look_up_data_12 ? _booth_data_0_T_1 : _booth_data_12_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_12_T_11 = 3'h5 == look_up_data_12 ? {{1'd0}, x_fu} : _booth_data_12_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_12_T_13 = 3'h6 == look_up_data_12 ? {{1'd0}, x_fu} : _booth_data_12_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_12_T_15 = 3'h7 == look_up_data_12 ? 133'h0 : _booth_data_12_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_12_T_17 = {1'h0,_booth_data_12_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [90:0] _GEN_11 = {_booth_data_12_T_17, 24'h0}; // @[hard_cal.scala 285:19]
  wire [97:0] _booth_data_12_T_18 = {{7'd0}, _GEN_11}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_13 = {regs_1[27],regs_1[26],regs_1[25]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_13_T_3 = 3'h1 == look_up_data_13 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_13_T_5 = 3'h2 == look_up_data_13 ? regs_0 : _booth_data_13_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_13_T_7 = 3'h3 == look_up_data_13 ? _booth_data_0_T : {{1'd0}, _booth_data_13_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_13_T_9 = 3'h4 == look_up_data_13 ? _booth_data_0_T_1 : _booth_data_13_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_13_T_11 = 3'h5 == look_up_data_13 ? {{1'd0}, x_fu} : _booth_data_13_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_13_T_13 = 3'h6 == look_up_data_13 ? {{1'd0}, x_fu} : _booth_data_13_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_13_T_15 = 3'h7 == look_up_data_13 ? 133'h0 : _booth_data_13_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_13_T_17 = {1'h0,_booth_data_13_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [92:0] _GEN_12 = {_booth_data_13_T_17, 26'h0}; // @[hard_cal.scala 285:19]
  wire [97:0] _booth_data_13_T_18 = {{5'd0}, _GEN_12}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_14 = {regs_1[29],regs_1[28],regs_1[27]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_14_T_3 = 3'h1 == look_up_data_14 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_14_T_5 = 3'h2 == look_up_data_14 ? regs_0 : _booth_data_14_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_14_T_7 = 3'h3 == look_up_data_14 ? _booth_data_0_T : {{1'd0}, _booth_data_14_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_14_T_9 = 3'h4 == look_up_data_14 ? _booth_data_0_T_1 : _booth_data_14_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_14_T_11 = 3'h5 == look_up_data_14 ? {{1'd0}, x_fu} : _booth_data_14_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_14_T_13 = 3'h6 == look_up_data_14 ? {{1'd0}, x_fu} : _booth_data_14_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_14_T_15 = 3'h7 == look_up_data_14 ? 133'h0 : _booth_data_14_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_14_T_17 = {1'h0,_booth_data_14_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [94:0] _GEN_13 = {_booth_data_14_T_17, 28'h0}; // @[hard_cal.scala 285:19]
  wire [97:0] _booth_data_14_T_18 = {{3'd0}, _GEN_13}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_15 = {regs_1[31],regs_1[30],regs_1[29]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_15_T_3 = 3'h1 == look_up_data_15 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_15_T_5 = 3'h2 == look_up_data_15 ? regs_0 : _booth_data_15_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_15_T_7 = 3'h3 == look_up_data_15 ? _booth_data_0_T : {{1'd0}, _booth_data_15_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_15_T_9 = 3'h4 == look_up_data_15 ? _booth_data_0_T_1 : _booth_data_15_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_15_T_11 = 3'h5 == look_up_data_15 ? {{1'd0}, x_fu} : _booth_data_15_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_15_T_13 = 3'h6 == look_up_data_15 ? {{1'd0}, x_fu} : _booth_data_15_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_15_T_15 = 3'h7 == look_up_data_15 ? 133'h0 : _booth_data_15_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_15_T_17 = {1'h0,_booth_data_15_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [96:0] _GEN_14 = {_booth_data_15_T_17, 30'h0}; // @[hard_cal.scala 285:19]
  wire [97:0] _booth_data_15_T_18 = {{1'd0}, _GEN_14}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_16 = {regs_1[33],regs_1[32],regs_1[31]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_16_T_3 = 3'h1 == look_up_data_16 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_16_T_5 = 3'h2 == look_up_data_16 ? regs_0 : _booth_data_16_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_16_T_7 = 3'h3 == look_up_data_16 ? _booth_data_0_T : {{1'd0}, _booth_data_16_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_16_T_9 = 3'h4 == look_up_data_16 ? _booth_data_0_T_1 : _booth_data_16_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_16_T_11 = 3'h5 == look_up_data_16 ? {{1'd0}, x_fu} : _booth_data_16_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_16_T_13 = 3'h6 == look_up_data_16 ? {{1'd0}, x_fu} : _booth_data_16_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_16_T_15 = 3'h7 == look_up_data_16 ? 133'h0 : _booth_data_16_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_16_T_17 = {1'h0,_booth_data_16_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [98:0] _GEN_15 = {_booth_data_16_T_17, 32'h0}; // @[hard_cal.scala 285:19]
  wire [129:0] _booth_data_16_T_18 = {{31'd0}, _GEN_15}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_17 = {regs_1[35],regs_1[34],regs_1[33]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_17_T_3 = 3'h1 == look_up_data_17 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_17_T_5 = 3'h2 == look_up_data_17 ? regs_0 : _booth_data_17_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_17_T_7 = 3'h3 == look_up_data_17 ? _booth_data_0_T : {{1'd0}, _booth_data_17_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_17_T_9 = 3'h4 == look_up_data_17 ? _booth_data_0_T_1 : _booth_data_17_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_17_T_11 = 3'h5 == look_up_data_17 ? {{1'd0}, x_fu} : _booth_data_17_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_17_T_13 = 3'h6 == look_up_data_17 ? {{1'd0}, x_fu} : _booth_data_17_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_17_T_15 = 3'h7 == look_up_data_17 ? 133'h0 : _booth_data_17_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_17_T_17 = {1'h0,_booth_data_17_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [100:0] _GEN_16 = {_booth_data_17_T_17, 34'h0}; // @[hard_cal.scala 285:19]
  wire [129:0] _booth_data_17_T_18 = {{29'd0}, _GEN_16}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_18 = {regs_1[37],regs_1[36],regs_1[35]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_18_T_3 = 3'h1 == look_up_data_18 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_18_T_5 = 3'h2 == look_up_data_18 ? regs_0 : _booth_data_18_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_18_T_7 = 3'h3 == look_up_data_18 ? _booth_data_0_T : {{1'd0}, _booth_data_18_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_18_T_9 = 3'h4 == look_up_data_18 ? _booth_data_0_T_1 : _booth_data_18_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_18_T_11 = 3'h5 == look_up_data_18 ? {{1'd0}, x_fu} : _booth_data_18_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_18_T_13 = 3'h6 == look_up_data_18 ? {{1'd0}, x_fu} : _booth_data_18_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_18_T_15 = 3'h7 == look_up_data_18 ? 133'h0 : _booth_data_18_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_18_T_17 = {1'h0,_booth_data_18_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [102:0] _GEN_17 = {_booth_data_18_T_17, 36'h0}; // @[hard_cal.scala 285:19]
  wire [129:0] _booth_data_18_T_18 = {{27'd0}, _GEN_17}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_19 = {regs_1[39],regs_1[38],regs_1[37]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_19_T_3 = 3'h1 == look_up_data_19 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_19_T_5 = 3'h2 == look_up_data_19 ? regs_0 : _booth_data_19_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_19_T_7 = 3'h3 == look_up_data_19 ? _booth_data_0_T : {{1'd0}, _booth_data_19_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_19_T_9 = 3'h4 == look_up_data_19 ? _booth_data_0_T_1 : _booth_data_19_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_19_T_11 = 3'h5 == look_up_data_19 ? {{1'd0}, x_fu} : _booth_data_19_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_19_T_13 = 3'h6 == look_up_data_19 ? {{1'd0}, x_fu} : _booth_data_19_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_19_T_15 = 3'h7 == look_up_data_19 ? 133'h0 : _booth_data_19_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_19_T_17 = {1'h0,_booth_data_19_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [104:0] _GEN_18 = {_booth_data_19_T_17, 38'h0}; // @[hard_cal.scala 285:19]
  wire [129:0] _booth_data_19_T_18 = {{25'd0}, _GEN_18}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_20 = {regs_1[41],regs_1[40],regs_1[39]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_20_T_3 = 3'h1 == look_up_data_20 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_20_T_5 = 3'h2 == look_up_data_20 ? regs_0 : _booth_data_20_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_20_T_7 = 3'h3 == look_up_data_20 ? _booth_data_0_T : {{1'd0}, _booth_data_20_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_20_T_9 = 3'h4 == look_up_data_20 ? _booth_data_0_T_1 : _booth_data_20_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_20_T_11 = 3'h5 == look_up_data_20 ? {{1'd0}, x_fu} : _booth_data_20_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_20_T_13 = 3'h6 == look_up_data_20 ? {{1'd0}, x_fu} : _booth_data_20_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_20_T_15 = 3'h7 == look_up_data_20 ? 133'h0 : _booth_data_20_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_20_T_17 = {1'h0,_booth_data_20_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [106:0] _GEN_19 = {_booth_data_20_T_17, 40'h0}; // @[hard_cal.scala 285:19]
  wire [129:0] _booth_data_20_T_18 = {{23'd0}, _GEN_19}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_21 = {regs_1[43],regs_1[42],regs_1[41]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_21_T_3 = 3'h1 == look_up_data_21 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_21_T_5 = 3'h2 == look_up_data_21 ? regs_0 : _booth_data_21_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_21_T_7 = 3'h3 == look_up_data_21 ? _booth_data_0_T : {{1'd0}, _booth_data_21_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_21_T_9 = 3'h4 == look_up_data_21 ? _booth_data_0_T_1 : _booth_data_21_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_21_T_11 = 3'h5 == look_up_data_21 ? {{1'd0}, x_fu} : _booth_data_21_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_21_T_13 = 3'h6 == look_up_data_21 ? {{1'd0}, x_fu} : _booth_data_21_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_21_T_15 = 3'h7 == look_up_data_21 ? 133'h0 : _booth_data_21_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_21_T_17 = {1'h0,_booth_data_21_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [108:0] _GEN_20 = {_booth_data_21_T_17, 42'h0}; // @[hard_cal.scala 285:19]
  wire [129:0] _booth_data_21_T_18 = {{21'd0}, _GEN_20}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_22 = {regs_1[45],regs_1[44],regs_1[43]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_22_T_3 = 3'h1 == look_up_data_22 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_22_T_5 = 3'h2 == look_up_data_22 ? regs_0 : _booth_data_22_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_22_T_7 = 3'h3 == look_up_data_22 ? _booth_data_0_T : {{1'd0}, _booth_data_22_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_22_T_9 = 3'h4 == look_up_data_22 ? _booth_data_0_T_1 : _booth_data_22_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_22_T_11 = 3'h5 == look_up_data_22 ? {{1'd0}, x_fu} : _booth_data_22_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_22_T_13 = 3'h6 == look_up_data_22 ? {{1'd0}, x_fu} : _booth_data_22_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_22_T_15 = 3'h7 == look_up_data_22 ? 133'h0 : _booth_data_22_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_22_T_17 = {1'h0,_booth_data_22_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [110:0] _GEN_21 = {_booth_data_22_T_17, 44'h0}; // @[hard_cal.scala 285:19]
  wire [129:0] _booth_data_22_T_18 = {{19'd0}, _GEN_21}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_23 = {regs_1[47],regs_1[46],regs_1[45]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_23_T_3 = 3'h1 == look_up_data_23 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_23_T_5 = 3'h2 == look_up_data_23 ? regs_0 : _booth_data_23_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_23_T_7 = 3'h3 == look_up_data_23 ? _booth_data_0_T : {{1'd0}, _booth_data_23_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_23_T_9 = 3'h4 == look_up_data_23 ? _booth_data_0_T_1 : _booth_data_23_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_23_T_11 = 3'h5 == look_up_data_23 ? {{1'd0}, x_fu} : _booth_data_23_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_23_T_13 = 3'h6 == look_up_data_23 ? {{1'd0}, x_fu} : _booth_data_23_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_23_T_15 = 3'h7 == look_up_data_23 ? 133'h0 : _booth_data_23_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_23_T_17 = {1'h0,_booth_data_23_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [112:0] _GEN_22 = {_booth_data_23_T_17, 46'h0}; // @[hard_cal.scala 285:19]
  wire [129:0] _booth_data_23_T_18 = {{17'd0}, _GEN_22}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_24 = {regs_1[49],regs_1[48],regs_1[47]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_24_T_3 = 3'h1 == look_up_data_24 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_24_T_5 = 3'h2 == look_up_data_24 ? regs_0 : _booth_data_24_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_24_T_7 = 3'h3 == look_up_data_24 ? _booth_data_0_T : {{1'd0}, _booth_data_24_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_24_T_9 = 3'h4 == look_up_data_24 ? _booth_data_0_T_1 : _booth_data_24_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_24_T_11 = 3'h5 == look_up_data_24 ? {{1'd0}, x_fu} : _booth_data_24_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_24_T_13 = 3'h6 == look_up_data_24 ? {{1'd0}, x_fu} : _booth_data_24_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_24_T_15 = 3'h7 == look_up_data_24 ? 133'h0 : _booth_data_24_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_24_T_17 = {1'h0,_booth_data_24_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [114:0] _GEN_23 = {_booth_data_24_T_17, 48'h0}; // @[hard_cal.scala 285:19]
  wire [129:0] _booth_data_24_T_18 = {{15'd0}, _GEN_23}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_25 = {regs_1[51],regs_1[50],regs_1[49]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_25_T_3 = 3'h1 == look_up_data_25 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_25_T_5 = 3'h2 == look_up_data_25 ? regs_0 : _booth_data_25_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_25_T_7 = 3'h3 == look_up_data_25 ? _booth_data_0_T : {{1'd0}, _booth_data_25_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_25_T_9 = 3'h4 == look_up_data_25 ? _booth_data_0_T_1 : _booth_data_25_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_25_T_11 = 3'h5 == look_up_data_25 ? {{1'd0}, x_fu} : _booth_data_25_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_25_T_13 = 3'h6 == look_up_data_25 ? {{1'd0}, x_fu} : _booth_data_25_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_25_T_15 = 3'h7 == look_up_data_25 ? 133'h0 : _booth_data_25_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_25_T_17 = {1'h0,_booth_data_25_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [116:0] _GEN_24 = {_booth_data_25_T_17, 50'h0}; // @[hard_cal.scala 285:19]
  wire [129:0] _booth_data_25_T_18 = {{13'd0}, _GEN_24}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_26 = {regs_1[53],regs_1[52],regs_1[51]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_26_T_3 = 3'h1 == look_up_data_26 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_26_T_5 = 3'h2 == look_up_data_26 ? regs_0 : _booth_data_26_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_26_T_7 = 3'h3 == look_up_data_26 ? _booth_data_0_T : {{1'd0}, _booth_data_26_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_26_T_9 = 3'h4 == look_up_data_26 ? _booth_data_0_T_1 : _booth_data_26_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_26_T_11 = 3'h5 == look_up_data_26 ? {{1'd0}, x_fu} : _booth_data_26_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_26_T_13 = 3'h6 == look_up_data_26 ? {{1'd0}, x_fu} : _booth_data_26_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_26_T_15 = 3'h7 == look_up_data_26 ? 133'h0 : _booth_data_26_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_26_T_17 = {1'h0,_booth_data_26_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [118:0] _GEN_25 = {_booth_data_26_T_17, 52'h0}; // @[hard_cal.scala 285:19]
  wire [129:0] _booth_data_26_T_18 = {{11'd0}, _GEN_25}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_27 = {regs_1[55],regs_1[54],regs_1[53]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_27_T_3 = 3'h1 == look_up_data_27 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_27_T_5 = 3'h2 == look_up_data_27 ? regs_0 : _booth_data_27_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_27_T_7 = 3'h3 == look_up_data_27 ? _booth_data_0_T : {{1'd0}, _booth_data_27_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_27_T_9 = 3'h4 == look_up_data_27 ? _booth_data_0_T_1 : _booth_data_27_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_27_T_11 = 3'h5 == look_up_data_27 ? {{1'd0}, x_fu} : _booth_data_27_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_27_T_13 = 3'h6 == look_up_data_27 ? {{1'd0}, x_fu} : _booth_data_27_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_27_T_15 = 3'h7 == look_up_data_27 ? 133'h0 : _booth_data_27_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_27_T_17 = {1'h0,_booth_data_27_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [120:0] _GEN_26 = {_booth_data_27_T_17, 54'h0}; // @[hard_cal.scala 285:19]
  wire [129:0] _booth_data_27_T_18 = {{9'd0}, _GEN_26}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_28 = {regs_1[57],regs_1[56],regs_1[55]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_28_T_3 = 3'h1 == look_up_data_28 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_28_T_5 = 3'h2 == look_up_data_28 ? regs_0 : _booth_data_28_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_28_T_7 = 3'h3 == look_up_data_28 ? _booth_data_0_T : {{1'd0}, _booth_data_28_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_28_T_9 = 3'h4 == look_up_data_28 ? _booth_data_0_T_1 : _booth_data_28_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_28_T_11 = 3'h5 == look_up_data_28 ? {{1'd0}, x_fu} : _booth_data_28_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_28_T_13 = 3'h6 == look_up_data_28 ? {{1'd0}, x_fu} : _booth_data_28_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_28_T_15 = 3'h7 == look_up_data_28 ? 133'h0 : _booth_data_28_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_28_T_17 = {1'h0,_booth_data_28_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [122:0] _GEN_27 = {_booth_data_28_T_17, 56'h0}; // @[hard_cal.scala 285:19]
  wire [129:0] _booth_data_28_T_18 = {{7'd0}, _GEN_27}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_29 = {regs_1[59],regs_1[58],regs_1[57]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_29_T_3 = 3'h1 == look_up_data_29 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_29_T_5 = 3'h2 == look_up_data_29 ? regs_0 : _booth_data_29_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_29_T_7 = 3'h3 == look_up_data_29 ? _booth_data_0_T : {{1'd0}, _booth_data_29_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_29_T_9 = 3'h4 == look_up_data_29 ? _booth_data_0_T_1 : _booth_data_29_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_29_T_11 = 3'h5 == look_up_data_29 ? {{1'd0}, x_fu} : _booth_data_29_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_29_T_13 = 3'h6 == look_up_data_29 ? {{1'd0}, x_fu} : _booth_data_29_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_29_T_15 = 3'h7 == look_up_data_29 ? 133'h0 : _booth_data_29_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_29_T_17 = {1'h0,_booth_data_29_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [124:0] _GEN_28 = {_booth_data_29_T_17, 58'h0}; // @[hard_cal.scala 285:19]
  wire [129:0] _booth_data_29_T_18 = {{5'd0}, _GEN_28}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_30 = {regs_1[61],regs_1[60],regs_1[59]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_30_T_3 = 3'h1 == look_up_data_30 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_30_T_5 = 3'h2 == look_up_data_30 ? regs_0 : _booth_data_30_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_30_T_7 = 3'h3 == look_up_data_30 ? _booth_data_0_T : {{1'd0}, _booth_data_30_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_30_T_9 = 3'h4 == look_up_data_30 ? _booth_data_0_T_1 : _booth_data_30_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_30_T_11 = 3'h5 == look_up_data_30 ? {{1'd0}, x_fu} : _booth_data_30_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_30_T_13 = 3'h6 == look_up_data_30 ? {{1'd0}, x_fu} : _booth_data_30_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_30_T_15 = 3'h7 == look_up_data_30 ? 133'h0 : _booth_data_30_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_30_T_17 = {1'h0,_booth_data_30_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [126:0] _GEN_29 = {_booth_data_30_T_17, 60'h0}; // @[hard_cal.scala 285:19]
  wire [129:0] _booth_data_30_T_18 = {{3'd0}, _GEN_29}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_31 = {regs_1[63],regs_1[62],regs_1[61]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_31_T_3 = 3'h1 == look_up_data_31 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_31_T_5 = 3'h2 == look_up_data_31 ? regs_0 : _booth_data_31_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_31_T_7 = 3'h3 == look_up_data_31 ? _booth_data_0_T : {{1'd0}, _booth_data_31_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_31_T_9 = 3'h4 == look_up_data_31 ? _booth_data_0_T_1 : _booth_data_31_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_31_T_11 = 3'h5 == look_up_data_31 ? {{1'd0}, x_fu} : _booth_data_31_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_31_T_13 = 3'h6 == look_up_data_31 ? {{1'd0}, x_fu} : _booth_data_31_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_31_T_15 = 3'h7 == look_up_data_31 ? 133'h0 : _booth_data_31_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_31_T_17 = {1'h0,_booth_data_31_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [128:0] _GEN_30 = {_booth_data_31_T_17, 62'h0}; // @[hard_cal.scala 285:19]
  wire [129:0] _booth_data_31_T_18 = {{1'd0}, _GEN_30}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_32 = {regs_1[65],regs_1[64],regs_1[63]}; // @[Cat.scala 31:58]
  wire [131:0] _booth_data_32_T_3 = 3'h1 == look_up_data_32 ? regs_0 : 132'h0; // @[Mux.scala 81:58]
  wire [131:0] _booth_data_32_T_5 = 3'h2 == look_up_data_32 ? regs_0 : _booth_data_32_T_3; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_32_T_7 = 3'h3 == look_up_data_32 ? _booth_data_0_T : {{1'd0}, _booth_data_32_T_5}; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_32_T_9 = 3'h4 == look_up_data_32 ? _booth_data_0_T_1 : _booth_data_32_T_7; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_32_T_11 = 3'h5 == look_up_data_32 ? {{1'd0}, x_fu} : _booth_data_32_T_9; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_32_T_13 = 3'h6 == look_up_data_32 ? {{1'd0}, x_fu} : _booth_data_32_T_11; // @[Mux.scala 81:58]
  wire [132:0] _booth_data_32_T_15 = 3'h7 == look_up_data_32 ? 133'h0 : _booth_data_32_T_13; // @[Mux.scala 81:58]
  wire [66:0] _booth_data_32_T_17 = {1'h0,_booth_data_32_T_15[65:0]}; // @[Cat.scala 31:58]
  wire [130:0] _GEN_31 = {_booth_data_32_T_17, 64'h0}; // @[hard_cal.scala 285:19]
  wire [193:0] _booth_data_32_T_18 = {{63'd0}, _GEN_31}; // @[hard_cal.scala 285:19]
  wire [65:0] _x_fu_T_1 = ~io_data_0; // @[hard_cal.scala 290:53]
  wire [65:0] _x_fu_T_3 = _x_fu_T_1 + 66'h1; // @[hard_cal.scala 290:67]
  wire [3:0] _cal_start_T_2 = 4'h9 - 4'h1; // @[hard_cal.scala 297:112]
  wire [6:0] _GEN_32 = {{3'd0}, _cal_start_T_2}; // @[hard_cal.scala 297:78]
  wire  _cal_start_T_4 = counter == _GEN_32 ? 1'h0 : cal_start; // @[hard_cal.scala 297:69]
  wallace_adder cal_module ( // @[hard_cal.scala 295:28]
    .clock(cal_module_clock),
    .reset(cal_module_reset),
    .io_data_in_0(cal_module_io_data_in_0),
    .io_data_in_1(cal_module_io_data_in_1),
    .io_data_in_2(cal_module_io_data_in_2),
    .io_data_in_3(cal_module_io_data_in_3),
    .io_data_in_4(cal_module_io_data_in_4),
    .io_data_in_5(cal_module_io_data_in_5),
    .io_data_in_6(cal_module_io_data_in_6),
    .io_data_in_7(cal_module_io_data_in_7),
    .io_data_in_8(cal_module_io_data_in_8),
    .io_data_in_9(cal_module_io_data_in_9),
    .io_data_in_10(cal_module_io_data_in_10),
    .io_data_in_11(cal_module_io_data_in_11),
    .io_data_in_12(cal_module_io_data_in_12),
    .io_data_in_13(cal_module_io_data_in_13),
    .io_data_in_14(cal_module_io_data_in_14),
    .io_data_in_15(cal_module_io_data_in_15),
    .io_data_in_16(cal_module_io_data_in_16),
    .io_data_in_17(cal_module_io_data_in_17),
    .io_data_in_18(cal_module_io_data_in_18),
    .io_data_in_19(cal_module_io_data_in_19),
    .io_data_in_20(cal_module_io_data_in_20),
    .io_data_in_21(cal_module_io_data_in_21),
    .io_data_in_22(cal_module_io_data_in_22),
    .io_data_in_23(cal_module_io_data_in_23),
    .io_data_in_24(cal_module_io_data_in_24),
    .io_data_in_25(cal_module_io_data_in_25),
    .io_data_in_26(cal_module_io_data_in_26),
    .io_data_in_27(cal_module_io_data_in_27),
    .io_data_in_28(cal_module_io_data_in_28),
    .io_data_in_29(cal_module_io_data_in_29),
    .io_data_in_30(cal_module_io_data_in_30),
    .io_data_in_31(cal_module_io_data_in_31),
    .io_data_in_32(cal_module_io_data_in_32),
    .io_result(cal_module_io_result)
  );
  assign io_result_0 = cal_start ? cal_module_io_result[65:0] : result_reg[65:0]; // @[hard_cal.scala 303:24]
  assign io_result_1 = cal_start ? cal_module_io_result[131:66] : result_reg[131:66]; // @[hard_cal.scala 304:24]
  assign io_input_ready = ~cal_start; // @[hard_cal.scala 306:23]
  assign io_Output_valid = counter == _GEN_32; // @[hard_cal.scala 305:34]
  assign cal_module_clock = clock;
  assign cal_module_reset = reset;
  assign cal_module_io_data_in_0 = {{64'd0}, _booth_data_0_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_1 = {{62'd0}, _booth_data_1_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_2 = {{58'd0}, _booth_data_2_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_3 = {{58'd0}, _booth_data_3_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_4 = {{50'd0}, _booth_data_4_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_5 = {{50'd0}, _booth_data_5_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_6 = {{50'd0}, _booth_data_6_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_7 = {{50'd0}, _booth_data_7_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_8 = {{34'd0}, _booth_data_8_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_9 = {{34'd0}, _booth_data_9_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_10 = {{34'd0}, _booth_data_10_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_11 = {{34'd0}, _booth_data_11_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_12 = {{34'd0}, _booth_data_12_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_13 = {{34'd0}, _booth_data_13_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_14 = {{34'd0}, _booth_data_14_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_15 = {{34'd0}, _booth_data_15_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_16 = {{2'd0}, _booth_data_16_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_17 = {{2'd0}, _booth_data_17_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_18 = {{2'd0}, _booth_data_18_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_19 = {{2'd0}, _booth_data_19_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_20 = {{2'd0}, _booth_data_20_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_21 = {{2'd0}, _booth_data_21_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_22 = {{2'd0}, _booth_data_22_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_23 = {{2'd0}, _booth_data_23_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_24 = {{2'd0}, _booth_data_24_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_25 = {{2'd0}, _booth_data_25_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_26 = {{2'd0}, _booth_data_26_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_27 = {{2'd0}, _booth_data_27_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_28 = {{2'd0}, _booth_data_28_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_29 = {{2'd0}, _booth_data_29_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_30 = {{2'd0}, _booth_data_30_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_31 = {{2'd0}, _booth_data_31_T_18}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_32 = _booth_data_32_T_18[131:0]; // @[hard_cal.scala 263:26 275:27]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 289:19]
      regs_0 <= 132'h0;
    end else if (_signed_T) begin
      regs_0 <= {{66'd0}, io_data_0};
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 291:19]
      regs_1 <= 132'h0;
    end else if (_signed_T) begin
      regs_1 <= {{66'd0}, io_data_1};
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 259:19]
      counter <= 7'h0;
    end else if (cal_start) begin
      counter <= _counter_T_1;
    end else begin
      counter <= 7'h0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 297:21]
      cal_start <= 1'h0;
    end else begin
      cal_start <= _signed_T | _cal_start_T_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 302:22]
      result_reg <= 132'h0;
    end else if (cal_start) begin
      result_reg <= cal_module_io_result;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 290:18]
      x_fu <= 132'h0;
    end else if (_signed_T) begin
      x_fu <= {{66'd0}, _x_fu_T_3};
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {5{`RANDOM}};
  regs_0 = _RAND_0[131:0];
  _RAND_1 = {5{`RANDOM}};
  regs_1 = _RAND_1[131:0];
  _RAND_2 = {1{`RANDOM}};
  counter = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  cal_start = _RAND_3[0:0];
  _RAND_4 = {5{`RANDOM}};
  result_reg = _RAND_4[131:0];
  _RAND_5 = {5{`RANDOM}};
  x_fu = _RAND_5[131:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    regs_0 = 132'h0;
  end
  if (reset) begin
    regs_1 = 132'h0;
  end
  if (reset) begin
    counter = 7'h0;
  end
  if (reset) begin
    cal_start = 1'h0;
  end
  if (reset) begin
    result_reg = 132'h0;
  end
  if (reset) begin
    x_fu = 132'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module csa_31(
  input  [67:0] io_data_0,
  input  [67:0] io_data_1,
  input  [67:0] io_data_2,
  output [67:0] io_result_0,
  output [67:0] io_result_1
);
  wire [67:0] _io_result_0_T = io_data_0 ^ io_data_1; // @[hard_cal.scala 182:32]
  wire [67:0] _io_result_1_T = io_data_0 & io_data_1; // @[hard_cal.scala 183:37]
  wire [67:0] _io_result_1_T_1 = io_data_1 & io_data_2; // @[hard_cal.scala 183:65]
  wire [67:0] _io_result_1_T_2 = _io_result_1_T | _io_result_1_T_1; // @[hard_cal.scala 183:51]
  wire [67:0] _io_result_1_T_3 = io_data_2 & io_data_0; // @[hard_cal.scala 183:93]
  wire [67:0] _io_result_1_T_4 = _io_result_1_T_2 | _io_result_1_T_3; // @[hard_cal.scala 183:79]
  wire [68:0] _io_result_1_T_5 = {_io_result_1_T_4,1'h0}; // @[Cat.scala 31:58]
  assign io_result_0 = _io_result_0_T ^ io_data_2; // @[hard_cal.scala 182:45]
  assign io_result_1 = _io_result_1_T_5[67:0]; // @[hard_cal.scala 183:18]
endmodule
module wallace_adder_1(
  input         clock,
  input         reset,
  input  [67:0] io_data_in_0,
  input  [67:0] io_data_in_1,
  input  [67:0] io_data_in_2,
  input  [67:0] io_data_in_3,
  input  [67:0] io_data_in_4,
  input  [67:0] io_data_in_5,
  input  [67:0] io_data_in_6,
  input  [67:0] io_data_in_7,
  input  [67:0] io_data_in_8,
  input  [67:0] io_data_in_9,
  input  [67:0] io_data_in_10,
  input  [67:0] io_data_in_11,
  input  [67:0] io_data_in_12,
  input  [67:0] io_data_in_13,
  input  [67:0] io_data_in_14,
  input  [67:0] io_data_in_15,
  input  [67:0] io_data_in_16,
  output [67:0] io_result
);
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [95:0] _RAND_2;
  reg [95:0] _RAND_3;
  reg [95:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [95:0] _RAND_6;
  reg [95:0] _RAND_7;
  reg [95:0] _RAND_8;
  reg [95:0] _RAND_9;
  reg [95:0] _RAND_10;
  reg [95:0] _RAND_11;
  reg [95:0] _RAND_12;
  reg [95:0] _RAND_13;
  reg [95:0] _RAND_14;
  reg [95:0] _RAND_15;
  reg [95:0] _RAND_16;
  reg [95:0] _RAND_17;
  reg [95:0] _RAND_18;
  reg [95:0] _RAND_19;
  reg [95:0] _RAND_20;
  reg [95:0] _RAND_21;
  reg [95:0] _RAND_22;
  reg [95:0] _RAND_23;
  reg [95:0] _RAND_24;
  reg [95:0] _RAND_25;
  reg [95:0] _RAND_26;
  reg [95:0] _RAND_27;
  reg [95:0] _RAND_28;
  reg [95:0] _RAND_29;
  reg [95:0] _RAND_30;
  reg [95:0] _RAND_31;
  reg [95:0] _RAND_32;
  reg [95:0] _RAND_33;
  reg [95:0] _RAND_34;
`endif // RANDOMIZE_REG_INIT
  wire [67:0] csa_io_data_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_io_data_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_io_data_2; // @[hard_cal.scala 204:61]
  wire [67:0] csa_io_result_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_io_result_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_1_io_data_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_1_io_data_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_1_io_data_2; // @[hard_cal.scala 204:61]
  wire [67:0] csa_1_io_result_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_1_io_result_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_2_io_data_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_2_io_data_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_2_io_data_2; // @[hard_cal.scala 204:61]
  wire [67:0] csa_2_io_result_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_2_io_result_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_3_io_data_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_3_io_data_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_3_io_data_2; // @[hard_cal.scala 204:61]
  wire [67:0] csa_3_io_result_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_3_io_result_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_4_io_data_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_4_io_data_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_4_io_data_2; // @[hard_cal.scala 204:61]
  wire [67:0] csa_4_io_result_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_4_io_result_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_5_io_data_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_5_io_data_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_5_io_data_2; // @[hard_cal.scala 204:61]
  wire [67:0] csa_5_io_result_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_5_io_result_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_6_io_data_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_6_io_data_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_6_io_data_2; // @[hard_cal.scala 204:61]
  wire [67:0] csa_6_io_result_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_6_io_result_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_7_io_data_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_7_io_data_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_7_io_data_2; // @[hard_cal.scala 204:61]
  wire [67:0] csa_7_io_result_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_7_io_result_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_8_io_data_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_8_io_data_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_8_io_data_2; // @[hard_cal.scala 204:61]
  wire [67:0] csa_8_io_result_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_8_io_result_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_9_io_data_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_9_io_data_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_9_io_data_2; // @[hard_cal.scala 204:61]
  wire [67:0] csa_9_io_result_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_9_io_result_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_10_io_data_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_10_io_data_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_10_io_data_2; // @[hard_cal.scala 204:61]
  wire [67:0] csa_10_io_result_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_10_io_result_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_11_io_data_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_11_io_data_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_11_io_data_2; // @[hard_cal.scala 204:61]
  wire [67:0] csa_11_io_result_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_11_io_result_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_12_io_data_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_12_io_data_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_12_io_data_2; // @[hard_cal.scala 204:61]
  wire [67:0] csa_12_io_result_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_12_io_result_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_13_io_data_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_13_io_data_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_13_io_data_2; // @[hard_cal.scala 204:61]
  wire [67:0] csa_13_io_result_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_13_io_result_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_14_io_data_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_14_io_data_1; // @[hard_cal.scala 204:61]
  wire [67:0] csa_14_io_data_2; // @[hard_cal.scala 204:61]
  wire [67:0] csa_14_io_result_0; // @[hard_cal.scala 204:61]
  wire [67:0] csa_14_io_result_1; // @[hard_cal.scala 204:61]
  reg [67:0] vec_data_out_data_reg__0; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg__1; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg__2; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg__3; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg__4; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg__5; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg__6; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg__7; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg__8; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg__9; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg__10; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg__11; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_1_0; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_1_1; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_1_2; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_1_3; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_1_4; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_1_5; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_1_6; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_1_7; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_2_0; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_2_1; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_2_2; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_2_3; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_2_4; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_2_5; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_3_0; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_3_1; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_3_2; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_3_3; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_4_0; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_4_1; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_out_data_reg_4_2; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_0; // @[hard_cal.scala 220:39]
  reg [67:0] vec_data_1; // @[hard_cal.scala 220:39]
  csa_31 csa ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_io_data_0),
    .io_data_1(csa_io_data_1),
    .io_data_2(csa_io_data_2),
    .io_result_0(csa_io_result_0),
    .io_result_1(csa_io_result_1)
  );
  csa_31 csa_1 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_1_io_data_0),
    .io_data_1(csa_1_io_data_1),
    .io_data_2(csa_1_io_data_2),
    .io_result_0(csa_1_io_result_0),
    .io_result_1(csa_1_io_result_1)
  );
  csa_31 csa_2 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_2_io_data_0),
    .io_data_1(csa_2_io_data_1),
    .io_data_2(csa_2_io_data_2),
    .io_result_0(csa_2_io_result_0),
    .io_result_1(csa_2_io_result_1)
  );
  csa_31 csa_3 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_3_io_data_0),
    .io_data_1(csa_3_io_data_1),
    .io_data_2(csa_3_io_data_2),
    .io_result_0(csa_3_io_result_0),
    .io_result_1(csa_3_io_result_1)
  );
  csa_31 csa_4 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_4_io_data_0),
    .io_data_1(csa_4_io_data_1),
    .io_data_2(csa_4_io_data_2),
    .io_result_0(csa_4_io_result_0),
    .io_result_1(csa_4_io_result_1)
  );
  csa_31 csa_5 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_5_io_data_0),
    .io_data_1(csa_5_io_data_1),
    .io_data_2(csa_5_io_data_2),
    .io_result_0(csa_5_io_result_0),
    .io_result_1(csa_5_io_result_1)
  );
  csa_31 csa_6 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_6_io_data_0),
    .io_data_1(csa_6_io_data_1),
    .io_data_2(csa_6_io_data_2),
    .io_result_0(csa_6_io_result_0),
    .io_result_1(csa_6_io_result_1)
  );
  csa_31 csa_7 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_7_io_data_0),
    .io_data_1(csa_7_io_data_1),
    .io_data_2(csa_7_io_data_2),
    .io_result_0(csa_7_io_result_0),
    .io_result_1(csa_7_io_result_1)
  );
  csa_31 csa_8 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_8_io_data_0),
    .io_data_1(csa_8_io_data_1),
    .io_data_2(csa_8_io_data_2),
    .io_result_0(csa_8_io_result_0),
    .io_result_1(csa_8_io_result_1)
  );
  csa_31 csa_9 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_9_io_data_0),
    .io_data_1(csa_9_io_data_1),
    .io_data_2(csa_9_io_data_2),
    .io_result_0(csa_9_io_result_0),
    .io_result_1(csa_9_io_result_1)
  );
  csa_31 csa_10 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_10_io_data_0),
    .io_data_1(csa_10_io_data_1),
    .io_data_2(csa_10_io_data_2),
    .io_result_0(csa_10_io_result_0),
    .io_result_1(csa_10_io_result_1)
  );
  csa_31 csa_11 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_11_io_data_0),
    .io_data_1(csa_11_io_data_1),
    .io_data_2(csa_11_io_data_2),
    .io_result_0(csa_11_io_result_0),
    .io_result_1(csa_11_io_result_1)
  );
  csa_31 csa_12 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_12_io_data_0),
    .io_data_1(csa_12_io_data_1),
    .io_data_2(csa_12_io_data_2),
    .io_result_0(csa_12_io_result_0),
    .io_result_1(csa_12_io_result_1)
  );
  csa_31 csa_13 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_13_io_data_0),
    .io_data_1(csa_13_io_data_1),
    .io_data_2(csa_13_io_data_2),
    .io_result_0(csa_13_io_result_0),
    .io_result_1(csa_13_io_result_1)
  );
  csa_31 csa_14 ( // @[hard_cal.scala 204:61]
    .io_data_0(csa_14_io_data_0),
    .io_data_1(csa_14_io_data_1),
    .io_data_2(csa_14_io_data_2),
    .io_result_0(csa_14_io_result_0),
    .io_result_1(csa_14_io_result_1)
  );
  assign io_result = vec_data_0 + vec_data_1; // @[hard_cal.scala 231:30]
  assign csa_io_data_0 = io_data_in_0; // @[hard_cal.scala 204:36 208:58]
  assign csa_io_data_1 = io_data_in_1; // @[hard_cal.scala 204:36 208:58]
  assign csa_io_data_2 = io_data_in_2; // @[hard_cal.scala 204:36 208:58]
  assign csa_1_io_data_0 = io_data_in_3; // @[hard_cal.scala 204:36 208:58]
  assign csa_1_io_data_1 = io_data_in_4; // @[hard_cal.scala 204:36 208:58]
  assign csa_1_io_data_2 = io_data_in_5; // @[hard_cal.scala 204:36 208:58]
  assign csa_2_io_data_0 = io_data_in_6; // @[hard_cal.scala 204:36 208:58]
  assign csa_2_io_data_1 = io_data_in_7; // @[hard_cal.scala 204:36 208:58]
  assign csa_2_io_data_2 = io_data_in_8; // @[hard_cal.scala 204:36 208:58]
  assign csa_3_io_data_0 = io_data_in_9; // @[hard_cal.scala 204:36 208:58]
  assign csa_3_io_data_1 = io_data_in_10; // @[hard_cal.scala 204:36 208:58]
  assign csa_3_io_data_2 = io_data_in_11; // @[hard_cal.scala 204:36 208:58]
  assign csa_4_io_data_0 = io_data_in_12; // @[hard_cal.scala 204:36 208:58]
  assign csa_4_io_data_1 = io_data_in_13; // @[hard_cal.scala 204:36 208:58]
  assign csa_4_io_data_2 = io_data_in_14; // @[hard_cal.scala 204:36 208:58]
  assign csa_5_io_data_0 = vec_data_out_data_reg__0; // @[hard_cal.scala 204:36 208:58]
  assign csa_5_io_data_1 = vec_data_out_data_reg__1; // @[hard_cal.scala 204:36 208:58]
  assign csa_5_io_data_2 = vec_data_out_data_reg__2; // @[hard_cal.scala 204:36 208:58]
  assign csa_6_io_data_0 = vec_data_out_data_reg__3; // @[hard_cal.scala 204:36 208:58]
  assign csa_6_io_data_1 = vec_data_out_data_reg__4; // @[hard_cal.scala 204:36 208:58]
  assign csa_6_io_data_2 = vec_data_out_data_reg__5; // @[hard_cal.scala 204:36 208:58]
  assign csa_7_io_data_0 = vec_data_out_data_reg__6; // @[hard_cal.scala 204:36 208:58]
  assign csa_7_io_data_1 = vec_data_out_data_reg__7; // @[hard_cal.scala 204:36 208:58]
  assign csa_7_io_data_2 = vec_data_out_data_reg__8; // @[hard_cal.scala 204:36 208:58]
  assign csa_8_io_data_0 = vec_data_out_data_reg__9; // @[hard_cal.scala 204:36 208:58]
  assign csa_8_io_data_1 = vec_data_out_data_reg__10; // @[hard_cal.scala 204:36 208:58]
  assign csa_8_io_data_2 = vec_data_out_data_reg__11; // @[hard_cal.scala 204:36 208:58]
  assign csa_9_io_data_0 = vec_data_out_data_reg_1_0; // @[hard_cal.scala 204:36 208:58]
  assign csa_9_io_data_1 = vec_data_out_data_reg_1_1; // @[hard_cal.scala 204:36 208:58]
  assign csa_9_io_data_2 = vec_data_out_data_reg_1_2; // @[hard_cal.scala 204:36 208:58]
  assign csa_10_io_data_0 = vec_data_out_data_reg_1_3; // @[hard_cal.scala 204:36 208:58]
  assign csa_10_io_data_1 = vec_data_out_data_reg_1_4; // @[hard_cal.scala 204:36 208:58]
  assign csa_10_io_data_2 = vec_data_out_data_reg_1_5; // @[hard_cal.scala 204:36 208:58]
  assign csa_11_io_data_0 = vec_data_out_data_reg_2_0; // @[hard_cal.scala 204:36 208:58]
  assign csa_11_io_data_1 = vec_data_out_data_reg_2_1; // @[hard_cal.scala 204:36 208:58]
  assign csa_11_io_data_2 = vec_data_out_data_reg_2_2; // @[hard_cal.scala 204:36 208:58]
  assign csa_12_io_data_0 = vec_data_out_data_reg_2_3; // @[hard_cal.scala 204:36 208:58]
  assign csa_12_io_data_1 = vec_data_out_data_reg_2_4; // @[hard_cal.scala 204:36 208:58]
  assign csa_12_io_data_2 = vec_data_out_data_reg_2_5; // @[hard_cal.scala 204:36 208:58]
  assign csa_13_io_data_0 = vec_data_out_data_reg_3_0; // @[hard_cal.scala 204:36 208:58]
  assign csa_13_io_data_1 = vec_data_out_data_reg_3_1; // @[hard_cal.scala 204:36 208:58]
  assign csa_13_io_data_2 = vec_data_out_data_reg_3_2; // @[hard_cal.scala 204:36 208:58]
  assign csa_14_io_data_0 = vec_data_out_data_reg_4_0; // @[hard_cal.scala 204:36 208:58]
  assign csa_14_io_data_1 = vec_data_out_data_reg_4_1; // @[hard_cal.scala 204:36 208:58]
  assign csa_14_io_data_2 = vec_data_out_data_reg_4_2; // @[hard_cal.scala 204:36 208:58]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__0 <= 68'h0;
    end else begin
      vec_data_out_data_reg__0 <= csa_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__1 <= 68'h0;
    end else begin
      vec_data_out_data_reg__1 <= csa_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__2 <= 68'h0;
    end else begin
      vec_data_out_data_reg__2 <= csa_1_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__3 <= 68'h0;
    end else begin
      vec_data_out_data_reg__3 <= csa_1_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__4 <= 68'h0;
    end else begin
      vec_data_out_data_reg__4 <= csa_2_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__5 <= 68'h0;
    end else begin
      vec_data_out_data_reg__5 <= csa_2_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__6 <= 68'h0;
    end else begin
      vec_data_out_data_reg__6 <= csa_3_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__7 <= 68'h0;
    end else begin
      vec_data_out_data_reg__7 <= csa_3_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__8 <= 68'h0;
    end else begin
      vec_data_out_data_reg__8 <= csa_4_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg__9 <= 68'h0;
    end else begin
      vec_data_out_data_reg__9 <= csa_4_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 211:39 217:44]
      vec_data_out_data_reg__10 <= 68'h0;
    end else begin
      vec_data_out_data_reg__10 <= io_data_in_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 211:39 217:44]
      vec_data_out_data_reg__11 <= 68'h0;
    end else begin
      vec_data_out_data_reg__11 <= io_data_in_16;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_0 <= 68'h0;
    end else begin
      vec_data_out_data_reg_1_0 <= csa_5_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_1 <= 68'h0;
    end else begin
      vec_data_out_data_reg_1_1 <= csa_5_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_2 <= 68'h0;
    end else begin
      vec_data_out_data_reg_1_2 <= csa_6_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_3 <= 68'h0;
    end else begin
      vec_data_out_data_reg_1_3 <= csa_6_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_4 <= 68'h0;
    end else begin
      vec_data_out_data_reg_1_4 <= csa_7_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_5 <= 68'h0;
    end else begin
      vec_data_out_data_reg_1_5 <= csa_7_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_6 <= 68'h0;
    end else begin
      vec_data_out_data_reg_1_6 <= csa_8_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_1_7 <= 68'h0;
    end else begin
      vec_data_out_data_reg_1_7 <= csa_8_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_2_0 <= 68'h0;
    end else begin
      vec_data_out_data_reg_2_0 <= csa_9_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_2_1 <= 68'h0;
    end else begin
      vec_data_out_data_reg_2_1 <= csa_9_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_2_2 <= 68'h0;
    end else begin
      vec_data_out_data_reg_2_2 <= csa_10_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_2_3 <= 68'h0;
    end else begin
      vec_data_out_data_reg_2_3 <= csa_10_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 211:39 217:44]
      vec_data_out_data_reg_2_4 <= 68'h0;
    end else begin
      vec_data_out_data_reg_2_4 <= vec_data_out_data_reg_1_6;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 211:39 217:44]
      vec_data_out_data_reg_2_5 <= 68'h0;
    end else begin
      vec_data_out_data_reg_2_5 <= vec_data_out_data_reg_1_7;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_3_0 <= 68'h0;
    end else begin
      vec_data_out_data_reg_3_0 <= csa_11_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_3_1 <= 68'h0;
    end else begin
      vec_data_out_data_reg_3_1 <= csa_11_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_3_2 <= 68'h0;
    end else begin
      vec_data_out_data_reg_3_2 <= csa_12_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_3_3 <= 68'h0;
    end else begin
      vec_data_out_data_reg_3_3 <= csa_12_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_4_0 <= 68'h0;
    end else begin
      vec_data_out_data_reg_4_0 <= csa_13_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_out_data_reg_4_1 <= 68'h0;
    end else begin
      vec_data_out_data_reg_4_1 <= csa_13_io_result_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 211:39 217:44]
      vec_data_out_data_reg_4_2 <= 68'h0;
    end else begin
      vec_data_out_data_reg_4_2 <= vec_data_out_data_reg_3_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_0 <= 68'h0;
    end else begin
      vec_data_0 <= csa_14_io_result_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 204:{36,36}]
      vec_data_1 <= 68'h0;
    end else begin
      vec_data_1 <= csa_14_io_result_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  vec_data_out_data_reg__0 = _RAND_0[67:0];
  _RAND_1 = {3{`RANDOM}};
  vec_data_out_data_reg__1 = _RAND_1[67:0];
  _RAND_2 = {3{`RANDOM}};
  vec_data_out_data_reg__2 = _RAND_2[67:0];
  _RAND_3 = {3{`RANDOM}};
  vec_data_out_data_reg__3 = _RAND_3[67:0];
  _RAND_4 = {3{`RANDOM}};
  vec_data_out_data_reg__4 = _RAND_4[67:0];
  _RAND_5 = {3{`RANDOM}};
  vec_data_out_data_reg__5 = _RAND_5[67:0];
  _RAND_6 = {3{`RANDOM}};
  vec_data_out_data_reg__6 = _RAND_6[67:0];
  _RAND_7 = {3{`RANDOM}};
  vec_data_out_data_reg__7 = _RAND_7[67:0];
  _RAND_8 = {3{`RANDOM}};
  vec_data_out_data_reg__8 = _RAND_8[67:0];
  _RAND_9 = {3{`RANDOM}};
  vec_data_out_data_reg__9 = _RAND_9[67:0];
  _RAND_10 = {3{`RANDOM}};
  vec_data_out_data_reg__10 = _RAND_10[67:0];
  _RAND_11 = {3{`RANDOM}};
  vec_data_out_data_reg__11 = _RAND_11[67:0];
  _RAND_12 = {3{`RANDOM}};
  vec_data_out_data_reg_1_0 = _RAND_12[67:0];
  _RAND_13 = {3{`RANDOM}};
  vec_data_out_data_reg_1_1 = _RAND_13[67:0];
  _RAND_14 = {3{`RANDOM}};
  vec_data_out_data_reg_1_2 = _RAND_14[67:0];
  _RAND_15 = {3{`RANDOM}};
  vec_data_out_data_reg_1_3 = _RAND_15[67:0];
  _RAND_16 = {3{`RANDOM}};
  vec_data_out_data_reg_1_4 = _RAND_16[67:0];
  _RAND_17 = {3{`RANDOM}};
  vec_data_out_data_reg_1_5 = _RAND_17[67:0];
  _RAND_18 = {3{`RANDOM}};
  vec_data_out_data_reg_1_6 = _RAND_18[67:0];
  _RAND_19 = {3{`RANDOM}};
  vec_data_out_data_reg_1_7 = _RAND_19[67:0];
  _RAND_20 = {3{`RANDOM}};
  vec_data_out_data_reg_2_0 = _RAND_20[67:0];
  _RAND_21 = {3{`RANDOM}};
  vec_data_out_data_reg_2_1 = _RAND_21[67:0];
  _RAND_22 = {3{`RANDOM}};
  vec_data_out_data_reg_2_2 = _RAND_22[67:0];
  _RAND_23 = {3{`RANDOM}};
  vec_data_out_data_reg_2_3 = _RAND_23[67:0];
  _RAND_24 = {3{`RANDOM}};
  vec_data_out_data_reg_2_4 = _RAND_24[67:0];
  _RAND_25 = {3{`RANDOM}};
  vec_data_out_data_reg_2_5 = _RAND_25[67:0];
  _RAND_26 = {3{`RANDOM}};
  vec_data_out_data_reg_3_0 = _RAND_26[67:0];
  _RAND_27 = {3{`RANDOM}};
  vec_data_out_data_reg_3_1 = _RAND_27[67:0];
  _RAND_28 = {3{`RANDOM}};
  vec_data_out_data_reg_3_2 = _RAND_28[67:0];
  _RAND_29 = {3{`RANDOM}};
  vec_data_out_data_reg_3_3 = _RAND_29[67:0];
  _RAND_30 = {3{`RANDOM}};
  vec_data_out_data_reg_4_0 = _RAND_30[67:0];
  _RAND_31 = {3{`RANDOM}};
  vec_data_out_data_reg_4_1 = _RAND_31[67:0];
  _RAND_32 = {3{`RANDOM}};
  vec_data_out_data_reg_4_2 = _RAND_32[67:0];
  _RAND_33 = {3{`RANDOM}};
  vec_data_0 = _RAND_33[67:0];
  _RAND_34 = {3{`RANDOM}};
  vec_data_1 = _RAND_34[67:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    vec_data_out_data_reg__0 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__1 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__2 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__3 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__4 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__5 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__6 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__7 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__8 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__9 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__10 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg__11 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_0 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_1 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_2 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_3 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_4 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_5 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_6 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_1_7 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_2_0 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_2_1 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_2_2 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_2_3 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_2_4 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_2_5 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_3_0 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_3_1 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_3_2 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_3_3 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_4_0 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_4_1 = 68'h0;
  end
  if (reset) begin
    vec_data_out_data_reg_4_2 = 68'h0;
  end
  if (reset) begin
    vec_data_0 = 68'h0;
  end
  if (reset) begin
    vec_data_1 = 68'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module mul_hard_1(
  input         clock,
  input         reset,
  output [33:0] io_result_0,
  input  [33:0] io_data_0,
  input  [33:0] io_data_1,
  input         io_input_valid,
  output        io_input_ready,
  output        io_Output_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [95:0] _RAND_4;
  reg [95:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  wire  cal_module_clock; // @[hard_cal.scala 295:28]
  wire  cal_module_reset; // @[hard_cal.scala 295:28]
  wire [67:0] cal_module_io_data_in_0; // @[hard_cal.scala 295:28]
  wire [67:0] cal_module_io_data_in_1; // @[hard_cal.scala 295:28]
  wire [67:0] cal_module_io_data_in_2; // @[hard_cal.scala 295:28]
  wire [67:0] cal_module_io_data_in_3; // @[hard_cal.scala 295:28]
  wire [67:0] cal_module_io_data_in_4; // @[hard_cal.scala 295:28]
  wire [67:0] cal_module_io_data_in_5; // @[hard_cal.scala 295:28]
  wire [67:0] cal_module_io_data_in_6; // @[hard_cal.scala 295:28]
  wire [67:0] cal_module_io_data_in_7; // @[hard_cal.scala 295:28]
  wire [67:0] cal_module_io_data_in_8; // @[hard_cal.scala 295:28]
  wire [67:0] cal_module_io_data_in_9; // @[hard_cal.scala 295:28]
  wire [67:0] cal_module_io_data_in_10; // @[hard_cal.scala 295:28]
  wire [67:0] cal_module_io_data_in_11; // @[hard_cal.scala 295:28]
  wire [67:0] cal_module_io_data_in_12; // @[hard_cal.scala 295:28]
  wire [67:0] cal_module_io_data_in_13; // @[hard_cal.scala 295:28]
  wire [67:0] cal_module_io_data_in_14; // @[hard_cal.scala 295:28]
  wire [67:0] cal_module_io_data_in_15; // @[hard_cal.scala 295:28]
  wire [67:0] cal_module_io_data_in_16; // @[hard_cal.scala 295:28]
  wire [67:0] cal_module_io_result; // @[hard_cal.scala 295:28]
  reg [67:0] regs_0; // @[hard_cal.scala 254:23]
  reg [67:0] regs_1; // @[hard_cal.scala 254:23]
  reg [5:0] counter; // @[hard_cal.scala 256:26]
  reg  cal_start; // @[hard_cal.scala 257:28]
  wire [5:0] _counter_T_1 = counter + 6'h1; // @[hard_cal.scala 259:39]
  wire  _signed_T = io_input_valid & io_input_ready; // @[hard_cal.scala 260:35]
  reg [67:0] result_reg; // @[hard_cal.scala 261:29]
  reg [67:0] x_fu; // @[hard_cal.scala 264:23]
  wire [2:0] look_up_data = {regs_1[1],regs_1[0],1'h0}; // @[Cat.scala 31:58]
  wire [68:0] _booth_data_0_T = {regs_0, 1'h0}; // @[hard_cal.scala 279:38]
  wire [68:0] _booth_data_0_T_1 = {x_fu, 1'h0}; // @[hard_cal.scala 280:31]
  wire [67:0] _booth_data_0_T_3 = 3'h1 == look_up_data ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_0_T_5 = 3'h2 == look_up_data ? regs_0 : _booth_data_0_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_0_T_7 = 3'h3 == look_up_data ? _booth_data_0_T : {{1'd0}, _booth_data_0_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_0_T_9 = 3'h4 == look_up_data ? _booth_data_0_T_1 : _booth_data_0_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_0_T_11 = 3'h5 == look_up_data ? {{1'd0}, x_fu} : _booth_data_0_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_0_T_13 = 3'h6 == look_up_data ? {{1'd0}, x_fu} : _booth_data_0_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_0_T_15 = 3'h7 == look_up_data ? 69'h0 : _booth_data_0_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_0_lo_lo = {_booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15[33],
    _booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_0_lo = {_booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15
    [33],_booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15[33],booth_data_0_lo_lo}
    ; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_0_T_46 = {_booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15[33],
    _booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15[33],_booth_data_0_T_15[33],
    booth_data_0_lo_lo,booth_data_0_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_0_T_48 = {_booth_data_0_T_46,_booth_data_0_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [64:0] _booth_data_0_T_49 = {{1'd0}, _booth_data_0_T_48}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_1 = {regs_1[3],regs_1[2],regs_1[1]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_1_T_3 = 3'h1 == look_up_data_1 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_1_T_5 = 3'h2 == look_up_data_1 ? regs_0 : _booth_data_1_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_1_T_7 = 3'h3 == look_up_data_1 ? _booth_data_0_T : {{1'd0}, _booth_data_1_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_1_T_9 = 3'h4 == look_up_data_1 ? _booth_data_0_T_1 : _booth_data_1_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_1_T_11 = 3'h5 == look_up_data_1 ? {{1'd0}, x_fu} : _booth_data_1_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_1_T_13 = 3'h6 == look_up_data_1 ? {{1'd0}, x_fu} : _booth_data_1_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_1_T_15 = 3'h7 == look_up_data_1 ? 69'h0 : _booth_data_1_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_1_lo_lo = {_booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15[33],
    _booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_1_lo = {_booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15
    [33],_booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15[33],booth_data_1_lo_lo}
    ; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_1_T_46 = {_booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15[33],
    _booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15[33],_booth_data_1_T_15[33],
    booth_data_1_lo_lo,booth_data_1_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_1_T_48 = {_booth_data_1_T_46,_booth_data_1_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [65:0] _GEN_0 = {_booth_data_1_T_48, 2'h0}; // @[hard_cal.scala 285:19]
  wire [66:0] _booth_data_1_T_49 = {{1'd0}, _GEN_0}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_2 = {regs_1[5],regs_1[4],regs_1[3]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_2_T_3 = 3'h1 == look_up_data_2 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_2_T_5 = 3'h2 == look_up_data_2 ? regs_0 : _booth_data_2_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_2_T_7 = 3'h3 == look_up_data_2 ? _booth_data_0_T : {{1'd0}, _booth_data_2_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_2_T_9 = 3'h4 == look_up_data_2 ? _booth_data_0_T_1 : _booth_data_2_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_2_T_11 = 3'h5 == look_up_data_2 ? {{1'd0}, x_fu} : _booth_data_2_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_2_T_13 = 3'h6 == look_up_data_2 ? {{1'd0}, x_fu} : _booth_data_2_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_2_T_15 = 3'h7 == look_up_data_2 ? 69'h0 : _booth_data_2_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_2_lo_lo = {_booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15[33],
    _booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_2_lo = {_booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15
    [33],_booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15[33],booth_data_2_lo_lo}
    ; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_2_T_46 = {_booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15[33],
    _booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15[33],_booth_data_2_T_15[33],
    booth_data_2_lo_lo,booth_data_2_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_2_T_48 = {_booth_data_2_T_46,_booth_data_2_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [67:0] _GEN_1 = {_booth_data_2_T_48, 4'h0}; // @[hard_cal.scala 285:19]
  wire [70:0] _booth_data_2_T_49 = {{3'd0}, _GEN_1}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_3 = {regs_1[7],regs_1[6],regs_1[5]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_3_T_3 = 3'h1 == look_up_data_3 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_3_T_5 = 3'h2 == look_up_data_3 ? regs_0 : _booth_data_3_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_3_T_7 = 3'h3 == look_up_data_3 ? _booth_data_0_T : {{1'd0}, _booth_data_3_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_3_T_9 = 3'h4 == look_up_data_3 ? _booth_data_0_T_1 : _booth_data_3_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_3_T_11 = 3'h5 == look_up_data_3 ? {{1'd0}, x_fu} : _booth_data_3_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_3_T_13 = 3'h6 == look_up_data_3 ? {{1'd0}, x_fu} : _booth_data_3_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_3_T_15 = 3'h7 == look_up_data_3 ? 69'h0 : _booth_data_3_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_3_lo_lo = {_booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15[33],
    _booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_3_lo = {_booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15
    [33],_booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15[33],booth_data_3_lo_lo}
    ; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_3_T_46 = {_booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15[33],
    _booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15[33],_booth_data_3_T_15[33],
    booth_data_3_lo_lo,booth_data_3_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_3_T_48 = {_booth_data_3_T_46,_booth_data_3_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [69:0] _GEN_2 = {_booth_data_3_T_48, 6'h0}; // @[hard_cal.scala 285:19]
  wire [70:0] _booth_data_3_T_49 = {{1'd0}, _GEN_2}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_4 = {regs_1[9],regs_1[8],regs_1[7]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_4_T_3 = 3'h1 == look_up_data_4 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_4_T_5 = 3'h2 == look_up_data_4 ? regs_0 : _booth_data_4_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_4_T_7 = 3'h3 == look_up_data_4 ? _booth_data_0_T : {{1'd0}, _booth_data_4_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_4_T_9 = 3'h4 == look_up_data_4 ? _booth_data_0_T_1 : _booth_data_4_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_4_T_11 = 3'h5 == look_up_data_4 ? {{1'd0}, x_fu} : _booth_data_4_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_4_T_13 = 3'h6 == look_up_data_4 ? {{1'd0}, x_fu} : _booth_data_4_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_4_T_15 = 3'h7 == look_up_data_4 ? 69'h0 : _booth_data_4_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_4_lo_lo = {_booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15[33],
    _booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_4_lo = {_booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15
    [33],_booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15[33],booth_data_4_lo_lo}
    ; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_4_T_46 = {_booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15[33],
    _booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15[33],_booth_data_4_T_15[33],
    booth_data_4_lo_lo,booth_data_4_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_4_T_48 = {_booth_data_4_T_46,_booth_data_4_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [71:0] _GEN_3 = {_booth_data_4_T_48, 8'h0}; // @[hard_cal.scala 285:19]
  wire [78:0] _booth_data_4_T_49 = {{7'd0}, _GEN_3}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_5 = {regs_1[11],regs_1[10],regs_1[9]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_5_T_3 = 3'h1 == look_up_data_5 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_5_T_5 = 3'h2 == look_up_data_5 ? regs_0 : _booth_data_5_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_5_T_7 = 3'h3 == look_up_data_5 ? _booth_data_0_T : {{1'd0}, _booth_data_5_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_5_T_9 = 3'h4 == look_up_data_5 ? _booth_data_0_T_1 : _booth_data_5_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_5_T_11 = 3'h5 == look_up_data_5 ? {{1'd0}, x_fu} : _booth_data_5_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_5_T_13 = 3'h6 == look_up_data_5 ? {{1'd0}, x_fu} : _booth_data_5_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_5_T_15 = 3'h7 == look_up_data_5 ? 69'h0 : _booth_data_5_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_5_lo_lo = {_booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15[33],
    _booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_5_lo = {_booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15
    [33],_booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15[33],booth_data_5_lo_lo}
    ; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_5_T_46 = {_booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15[33],
    _booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15[33],_booth_data_5_T_15[33],
    booth_data_5_lo_lo,booth_data_5_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_5_T_48 = {_booth_data_5_T_46,_booth_data_5_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [73:0] _GEN_4 = {_booth_data_5_T_48, 10'h0}; // @[hard_cal.scala 285:19]
  wire [78:0] _booth_data_5_T_49 = {{5'd0}, _GEN_4}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_6 = {regs_1[13],regs_1[12],regs_1[11]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_6_T_3 = 3'h1 == look_up_data_6 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_6_T_5 = 3'h2 == look_up_data_6 ? regs_0 : _booth_data_6_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_6_T_7 = 3'h3 == look_up_data_6 ? _booth_data_0_T : {{1'd0}, _booth_data_6_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_6_T_9 = 3'h4 == look_up_data_6 ? _booth_data_0_T_1 : _booth_data_6_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_6_T_11 = 3'h5 == look_up_data_6 ? {{1'd0}, x_fu} : _booth_data_6_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_6_T_13 = 3'h6 == look_up_data_6 ? {{1'd0}, x_fu} : _booth_data_6_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_6_T_15 = 3'h7 == look_up_data_6 ? 69'h0 : _booth_data_6_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_6_lo_lo = {_booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15[33],
    _booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_6_lo = {_booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15
    [33],_booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15[33],booth_data_6_lo_lo}
    ; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_6_T_46 = {_booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15[33],
    _booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15[33],_booth_data_6_T_15[33],
    booth_data_6_lo_lo,booth_data_6_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_6_T_48 = {_booth_data_6_T_46,_booth_data_6_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [75:0] _GEN_5 = {_booth_data_6_T_48, 12'h0}; // @[hard_cal.scala 285:19]
  wire [78:0] _booth_data_6_T_49 = {{3'd0}, _GEN_5}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_7 = {regs_1[15],regs_1[14],regs_1[13]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_7_T_3 = 3'h1 == look_up_data_7 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_7_T_5 = 3'h2 == look_up_data_7 ? regs_0 : _booth_data_7_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_7_T_7 = 3'h3 == look_up_data_7 ? _booth_data_0_T : {{1'd0}, _booth_data_7_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_7_T_9 = 3'h4 == look_up_data_7 ? _booth_data_0_T_1 : _booth_data_7_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_7_T_11 = 3'h5 == look_up_data_7 ? {{1'd0}, x_fu} : _booth_data_7_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_7_T_13 = 3'h6 == look_up_data_7 ? {{1'd0}, x_fu} : _booth_data_7_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_7_T_15 = 3'h7 == look_up_data_7 ? 69'h0 : _booth_data_7_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_7_lo_lo = {_booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15[33],
    _booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_7_lo = {_booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15
    [33],_booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15[33],booth_data_7_lo_lo}
    ; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_7_T_46 = {_booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15[33],
    _booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15[33],_booth_data_7_T_15[33],
    booth_data_7_lo_lo,booth_data_7_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_7_T_48 = {_booth_data_7_T_46,_booth_data_7_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [77:0] _GEN_6 = {_booth_data_7_T_48, 14'h0}; // @[hard_cal.scala 285:19]
  wire [78:0] _booth_data_7_T_49 = {{1'd0}, _GEN_6}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_8 = {regs_1[17],regs_1[16],regs_1[15]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_8_T_3 = 3'h1 == look_up_data_8 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_8_T_5 = 3'h2 == look_up_data_8 ? regs_0 : _booth_data_8_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_8_T_7 = 3'h3 == look_up_data_8 ? _booth_data_0_T : {{1'd0}, _booth_data_8_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_8_T_9 = 3'h4 == look_up_data_8 ? _booth_data_0_T_1 : _booth_data_8_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_8_T_11 = 3'h5 == look_up_data_8 ? {{1'd0}, x_fu} : _booth_data_8_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_8_T_13 = 3'h6 == look_up_data_8 ? {{1'd0}, x_fu} : _booth_data_8_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_8_T_15 = 3'h7 == look_up_data_8 ? 69'h0 : _booth_data_8_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_8_lo_lo = {_booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15[33],
    _booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_8_lo = {_booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15
    [33],_booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15[33],booth_data_8_lo_lo}
    ; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_8_T_46 = {_booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15[33],
    _booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15[33],_booth_data_8_T_15[33],
    booth_data_8_lo_lo,booth_data_8_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_8_T_48 = {_booth_data_8_T_46,_booth_data_8_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [79:0] _GEN_7 = {_booth_data_8_T_48, 16'h0}; // @[hard_cal.scala 285:19]
  wire [94:0] _booth_data_8_T_49 = {{15'd0}, _GEN_7}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_9 = {regs_1[19],regs_1[18],regs_1[17]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_9_T_3 = 3'h1 == look_up_data_9 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_9_T_5 = 3'h2 == look_up_data_9 ? regs_0 : _booth_data_9_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_9_T_7 = 3'h3 == look_up_data_9 ? _booth_data_0_T : {{1'd0}, _booth_data_9_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_9_T_9 = 3'h4 == look_up_data_9 ? _booth_data_0_T_1 : _booth_data_9_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_9_T_11 = 3'h5 == look_up_data_9 ? {{1'd0}, x_fu} : _booth_data_9_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_9_T_13 = 3'h6 == look_up_data_9 ? {{1'd0}, x_fu} : _booth_data_9_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_9_T_15 = 3'h7 == look_up_data_9 ? 69'h0 : _booth_data_9_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_9_lo_lo = {_booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15[33],
    _booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_9_lo = {_booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15
    [33],_booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15[33],booth_data_9_lo_lo}
    ; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_9_T_46 = {_booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15[33],
    _booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15[33],_booth_data_9_T_15[33],
    booth_data_9_lo_lo,booth_data_9_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_9_T_48 = {_booth_data_9_T_46,_booth_data_9_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [81:0] _GEN_8 = {_booth_data_9_T_48, 18'h0}; // @[hard_cal.scala 285:19]
  wire [94:0] _booth_data_9_T_49 = {{13'd0}, _GEN_8}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_10 = {regs_1[21],regs_1[20],regs_1[19]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_10_T_3 = 3'h1 == look_up_data_10 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_10_T_5 = 3'h2 == look_up_data_10 ? regs_0 : _booth_data_10_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_10_T_7 = 3'h3 == look_up_data_10 ? _booth_data_0_T : {{1'd0}, _booth_data_10_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_10_T_9 = 3'h4 == look_up_data_10 ? _booth_data_0_T_1 : _booth_data_10_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_10_T_11 = 3'h5 == look_up_data_10 ? {{1'd0}, x_fu} : _booth_data_10_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_10_T_13 = 3'h6 == look_up_data_10 ? {{1'd0}, x_fu} : _booth_data_10_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_10_T_15 = 3'h7 == look_up_data_10 ? 69'h0 : _booth_data_10_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_10_lo_lo = {_booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[33],
    _booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_10_lo = {_booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[33],
    _booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[
    33],booth_data_10_lo_lo}; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_10_T_46 = {_booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[33],
    _booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[33],_booth_data_10_T_15[
    33],booth_data_10_lo_lo,booth_data_10_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_10_T_48 = {_booth_data_10_T_46,_booth_data_10_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [83:0] _GEN_9 = {_booth_data_10_T_48, 20'h0}; // @[hard_cal.scala 285:19]
  wire [94:0] _booth_data_10_T_49 = {{11'd0}, _GEN_9}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_11 = {regs_1[23],regs_1[22],regs_1[21]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_11_T_3 = 3'h1 == look_up_data_11 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_11_T_5 = 3'h2 == look_up_data_11 ? regs_0 : _booth_data_11_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_11_T_7 = 3'h3 == look_up_data_11 ? _booth_data_0_T : {{1'd0}, _booth_data_11_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_11_T_9 = 3'h4 == look_up_data_11 ? _booth_data_0_T_1 : _booth_data_11_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_11_T_11 = 3'h5 == look_up_data_11 ? {{1'd0}, x_fu} : _booth_data_11_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_11_T_13 = 3'h6 == look_up_data_11 ? {{1'd0}, x_fu} : _booth_data_11_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_11_T_15 = 3'h7 == look_up_data_11 ? 69'h0 : _booth_data_11_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_11_lo_lo = {_booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[33],
    _booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_11_lo = {_booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[33],
    _booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[
    33],booth_data_11_lo_lo}; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_11_T_46 = {_booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[33],
    _booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[33],_booth_data_11_T_15[
    33],booth_data_11_lo_lo,booth_data_11_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_11_T_48 = {_booth_data_11_T_46,_booth_data_11_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [85:0] _GEN_10 = {_booth_data_11_T_48, 22'h0}; // @[hard_cal.scala 285:19]
  wire [94:0] _booth_data_11_T_49 = {{9'd0}, _GEN_10}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_12 = {regs_1[25],regs_1[24],regs_1[23]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_12_T_3 = 3'h1 == look_up_data_12 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_12_T_5 = 3'h2 == look_up_data_12 ? regs_0 : _booth_data_12_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_12_T_7 = 3'h3 == look_up_data_12 ? _booth_data_0_T : {{1'd0}, _booth_data_12_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_12_T_9 = 3'h4 == look_up_data_12 ? _booth_data_0_T_1 : _booth_data_12_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_12_T_11 = 3'h5 == look_up_data_12 ? {{1'd0}, x_fu} : _booth_data_12_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_12_T_13 = 3'h6 == look_up_data_12 ? {{1'd0}, x_fu} : _booth_data_12_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_12_T_15 = 3'h7 == look_up_data_12 ? 69'h0 : _booth_data_12_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_12_lo_lo = {_booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[33],
    _booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_12_lo = {_booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[33],
    _booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[
    33],booth_data_12_lo_lo}; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_12_T_46 = {_booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[33],
    _booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[33],_booth_data_12_T_15[
    33],booth_data_12_lo_lo,booth_data_12_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_12_T_48 = {_booth_data_12_T_46,_booth_data_12_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [87:0] _GEN_11 = {_booth_data_12_T_48, 24'h0}; // @[hard_cal.scala 285:19]
  wire [94:0] _booth_data_12_T_49 = {{7'd0}, _GEN_11}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_13 = {regs_1[27],regs_1[26],regs_1[25]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_13_T_3 = 3'h1 == look_up_data_13 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_13_T_5 = 3'h2 == look_up_data_13 ? regs_0 : _booth_data_13_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_13_T_7 = 3'h3 == look_up_data_13 ? _booth_data_0_T : {{1'd0}, _booth_data_13_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_13_T_9 = 3'h4 == look_up_data_13 ? _booth_data_0_T_1 : _booth_data_13_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_13_T_11 = 3'h5 == look_up_data_13 ? {{1'd0}, x_fu} : _booth_data_13_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_13_T_13 = 3'h6 == look_up_data_13 ? {{1'd0}, x_fu} : _booth_data_13_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_13_T_15 = 3'h7 == look_up_data_13 ? 69'h0 : _booth_data_13_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_13_lo_lo = {_booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[33],
    _booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_13_lo = {_booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[33],
    _booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[
    33],booth_data_13_lo_lo}; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_13_T_46 = {_booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[33],
    _booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[33],_booth_data_13_T_15[
    33],booth_data_13_lo_lo,booth_data_13_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_13_T_48 = {_booth_data_13_T_46,_booth_data_13_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [89:0] _GEN_12 = {_booth_data_13_T_48, 26'h0}; // @[hard_cal.scala 285:19]
  wire [94:0] _booth_data_13_T_49 = {{5'd0}, _GEN_12}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_14 = {regs_1[29],regs_1[28],regs_1[27]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_14_T_3 = 3'h1 == look_up_data_14 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_14_T_5 = 3'h2 == look_up_data_14 ? regs_0 : _booth_data_14_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_14_T_7 = 3'h3 == look_up_data_14 ? _booth_data_0_T : {{1'd0}, _booth_data_14_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_14_T_9 = 3'h4 == look_up_data_14 ? _booth_data_0_T_1 : _booth_data_14_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_14_T_11 = 3'h5 == look_up_data_14 ? {{1'd0}, x_fu} : _booth_data_14_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_14_T_13 = 3'h6 == look_up_data_14 ? {{1'd0}, x_fu} : _booth_data_14_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_14_T_15 = 3'h7 == look_up_data_14 ? 69'h0 : _booth_data_14_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_14_lo_lo = {_booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[33],
    _booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_14_lo = {_booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[33],
    _booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[
    33],booth_data_14_lo_lo}; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_14_T_46 = {_booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[33],
    _booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[33],_booth_data_14_T_15[
    33],booth_data_14_lo_lo,booth_data_14_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_14_T_48 = {_booth_data_14_T_46,_booth_data_14_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [91:0] _GEN_13 = {_booth_data_14_T_48, 28'h0}; // @[hard_cal.scala 285:19]
  wire [94:0] _booth_data_14_T_49 = {{3'd0}, _GEN_13}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_15 = {regs_1[31],regs_1[30],regs_1[29]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_15_T_3 = 3'h1 == look_up_data_15 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_15_T_5 = 3'h2 == look_up_data_15 ? regs_0 : _booth_data_15_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_15_T_7 = 3'h3 == look_up_data_15 ? _booth_data_0_T : {{1'd0}, _booth_data_15_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_15_T_9 = 3'h4 == look_up_data_15 ? _booth_data_0_T_1 : _booth_data_15_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_15_T_11 = 3'h5 == look_up_data_15 ? {{1'd0}, x_fu} : _booth_data_15_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_15_T_13 = 3'h6 == look_up_data_15 ? {{1'd0}, x_fu} : _booth_data_15_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_15_T_15 = 3'h7 == look_up_data_15 ? 69'h0 : _booth_data_15_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_15_lo_lo = {_booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[33],
    _booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_15_lo = {_booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[33],
    _booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[
    33],booth_data_15_lo_lo}; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_15_T_46 = {_booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[33],
    _booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[33],_booth_data_15_T_15[
    33],booth_data_15_lo_lo,booth_data_15_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_15_T_48 = {_booth_data_15_T_46,_booth_data_15_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [93:0] _GEN_14 = {_booth_data_15_T_48, 30'h0}; // @[hard_cal.scala 285:19]
  wire [94:0] _booth_data_15_T_49 = {{1'd0}, _GEN_14}; // @[hard_cal.scala 285:19]
  wire [2:0] look_up_data_16 = {regs_1[33],regs_1[32],regs_1[31]}; // @[Cat.scala 31:58]
  wire [67:0] _booth_data_16_T_3 = 3'h1 == look_up_data_16 ? regs_0 : 68'h0; // @[Mux.scala 81:58]
  wire [67:0] _booth_data_16_T_5 = 3'h2 == look_up_data_16 ? regs_0 : _booth_data_16_T_3; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_16_T_7 = 3'h3 == look_up_data_16 ? _booth_data_0_T : {{1'd0}, _booth_data_16_T_5}; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_16_T_9 = 3'h4 == look_up_data_16 ? _booth_data_0_T_1 : _booth_data_16_T_7; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_16_T_11 = 3'h5 == look_up_data_16 ? {{1'd0}, x_fu} : _booth_data_16_T_9; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_16_T_13 = 3'h6 == look_up_data_16 ? {{1'd0}, x_fu} : _booth_data_16_T_11; // @[Mux.scala 81:58]
  wire [68:0] _booth_data_16_T_15 = 3'h7 == look_up_data_16 ? 69'h0 : _booth_data_16_T_13; // @[Mux.scala 81:58]
  wire [6:0] booth_data_16_lo_lo = {_booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[33],
    _booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[33]}; // @[Cat.scala 31:58]
  wire [14:0] booth_data_16_lo = {_booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[33],
    _booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[
    33],booth_data_16_lo_lo}; // @[Cat.scala 31:58]
  wire [29:0] _booth_data_16_T_46 = {_booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[33],
    _booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[33],_booth_data_16_T_15[
    33],booth_data_16_lo_lo,booth_data_16_lo}; // @[Cat.scala 31:58]
  wire [63:0] _booth_data_16_T_48 = {_booth_data_16_T_46,_booth_data_16_T_15[33:0]}; // @[Cat.scala 31:58]
  wire [95:0] _GEN_15 = {_booth_data_16_T_48, 32'h0}; // @[hard_cal.scala 285:19]
  wire [126:0] _booth_data_16_T_49 = {{31'd0}, _GEN_15}; // @[hard_cal.scala 285:19]
  wire [33:0] _x_fu_T_1 = ~io_data_0; // @[hard_cal.scala 290:53]
  wire [33:0] _x_fu_T_3 = _x_fu_T_1 + 34'h1; // @[hard_cal.scala 290:67]
  wire [2:0] _cal_start_T_2 = 3'h7 - 3'h1; // @[hard_cal.scala 297:112]
  wire [5:0] _GEN_16 = {{3'd0}, _cal_start_T_2}; // @[hard_cal.scala 297:78]
  wire  _cal_start_T_4 = counter == _GEN_16 ? 1'h0 : cal_start; // @[hard_cal.scala 297:69]
  wallace_adder_1 cal_module ( // @[hard_cal.scala 295:28]
    .clock(cal_module_clock),
    .reset(cal_module_reset),
    .io_data_in_0(cal_module_io_data_in_0),
    .io_data_in_1(cal_module_io_data_in_1),
    .io_data_in_2(cal_module_io_data_in_2),
    .io_data_in_3(cal_module_io_data_in_3),
    .io_data_in_4(cal_module_io_data_in_4),
    .io_data_in_5(cal_module_io_data_in_5),
    .io_data_in_6(cal_module_io_data_in_6),
    .io_data_in_7(cal_module_io_data_in_7),
    .io_data_in_8(cal_module_io_data_in_8),
    .io_data_in_9(cal_module_io_data_in_9),
    .io_data_in_10(cal_module_io_data_in_10),
    .io_data_in_11(cal_module_io_data_in_11),
    .io_data_in_12(cal_module_io_data_in_12),
    .io_data_in_13(cal_module_io_data_in_13),
    .io_data_in_14(cal_module_io_data_in_14),
    .io_data_in_15(cal_module_io_data_in_15),
    .io_data_in_16(cal_module_io_data_in_16),
    .io_result(cal_module_io_result)
  );
  assign io_result_0 = cal_start ? cal_module_io_result[33:0] : result_reg[33:0]; // @[hard_cal.scala 303:24]
  assign io_input_ready = ~cal_start; // @[hard_cal.scala 306:23]
  assign io_Output_valid = counter == _GEN_16; // @[hard_cal.scala 305:34]
  assign cal_module_clock = clock;
  assign cal_module_reset = reset;
  assign cal_module_io_data_in_0 = {{3'd0}, _booth_data_0_T_49}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_1 = {{1'd0}, _booth_data_1_T_49}; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_2 = _booth_data_2_T_49[67:0]; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_3 = _booth_data_3_T_49[67:0]; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_4 = _booth_data_4_T_49[67:0]; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_5 = _booth_data_5_T_49[67:0]; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_6 = _booth_data_6_T_49[67:0]; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_7 = _booth_data_7_T_49[67:0]; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_8 = _booth_data_8_T_49[67:0]; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_9 = _booth_data_9_T_49[67:0]; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_10 = _booth_data_10_T_49[67:0]; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_11 = _booth_data_11_T_49[67:0]; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_12 = _booth_data_12_T_49[67:0]; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_13 = _booth_data_13_T_49[67:0]; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_14 = _booth_data_14_T_49[67:0]; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_15 = _booth_data_15_T_49[67:0]; // @[hard_cal.scala 263:26 275:27]
  assign cal_module_io_data_in_16 = _booth_data_16_T_49[67:0]; // @[hard_cal.scala 263:26 275:27]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 289:19]
      regs_0 <= 68'h0;
    end else if (_signed_T) begin
      regs_0 <= {{34'd0}, io_data_0};
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 291:19]
      regs_1 <= 68'h0;
    end else if (_signed_T) begin
      regs_1 <= {{34'd0}, io_data_1};
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 259:19]
      counter <= 6'h0;
    end else if (cal_start) begin
      counter <= _counter_T_1;
    end else begin
      counter <= 6'h0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 297:21]
      cal_start <= 1'h0;
    end else begin
      cal_start <= _signed_T | _cal_start_T_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 302:22]
      result_reg <= 68'h0;
    end else if (cal_start) begin
      result_reg <= cal_module_io_result;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 290:18]
      x_fu <= 68'h0;
    end else if (_signed_T) begin
      x_fu <= {{34'd0}, _x_fu_T_3};
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  regs_0 = _RAND_0[67:0];
  _RAND_1 = {3{`RANDOM}};
  regs_1 = _RAND_1[67:0];
  _RAND_2 = {1{`RANDOM}};
  counter = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  cal_start = _RAND_3[0:0];
  _RAND_4 = {3{`RANDOM}};
  result_reg = _RAND_4[67:0];
  _RAND_5 = {3{`RANDOM}};
  x_fu = _RAND_5[67:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    regs_0 = 68'h0;
  end
  if (reset) begin
    regs_1 = 68'h0;
  end
  if (reset) begin
    counter = 6'h0;
  end
  if (reset) begin
    cal_start = 1'h0;
  end
  if (reset) begin
    result_reg = 68'h0;
  end
  if (reset) begin
    x_fu = 68'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module div_simple(
  input         clock,
  input         reset,
  output [63:0] io_result_0,
  output [63:0] io_result_1,
  input  [63:0] io_data_0,
  input  [63:0] io_data_1,
  input         io_input_valid,
  output        io_input_ready,
  output        io_Output_valid,
  input         io_signed
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] regs_0; // @[hard_cal.scala 63:23]
  reg [127:0] regs_1; // @[hard_cal.scala 63:23]
  reg [6:0] counter; // @[hard_cal.scala 65:26]
  reg  cal_start; // @[hard_cal.scala 66:28]
  wire  _cal_start_T = io_input_valid & io_input_ready; // @[hard_cal.scala 67:37]
  wire  _cal_start_T_2 = counter == 7'h40 ? 1'h0 : cal_start; // @[hard_cal.scala 67:69]
  wire [6:0] _counter_T_1 = counter + 7'h1; // @[hard_cal.scala 68:39]
  reg [63:0] result_reg; // @[hard_cal.scala 70:29]
  wire [63:0] _data_in_0_T_2 = ~io_data_0; // @[hard_cal.scala 74:59]
  wire [63:0] _data_in_0_T_4 = _data_in_0_T_2 + 64'h1; // @[hard_cal.scala 74:76]
  wire [63:0] data_in_0 = io_signed & io_data_0[63] ? _data_in_0_T_4 : io_data_0; // @[hard_cal.scala 74:17]
  wire [63:0] _data_in_1_T_2 = ~io_data_1; // @[hard_cal.scala 74:59]
  wire [63:0] _data_in_1_T_4 = _data_in_1_T_2 + 64'h1; // @[hard_cal.scala 74:76]
  wire [63:0] data_in_1 = io_signed & io_data_1[63] ? _data_in_1_T_4 : io_data_1; // @[hard_cal.scala 74:17]
  wire [1:0] _T_2 = {io_data_0[63],io_data_1[63]}; // @[Cat.scala 31:58]
  wire  _T_6_1 = 2'h1 == _T_2 ? 1'h0 : 1'h1; // @[Mux.scala 81:58]
  wire  _T_8_0 = 2'h0 == _T_2 ? 1'h0 : 2'h1 == _T_2 | 2'h2 == _T_2; // @[Mux.scala 81:58]
  wire  _T_8_1 = 2'h0 == _T_2 ? 1'h0 : _T_6_1; // @[Mux.scala 81:58]
  wire  result_sign_0 = io_signed & _T_8_0; // @[hard_cal.scala 77:23]
  wire  result_sign_1 = io_signed & _T_8_1; // @[hard_cal.scala 77:23]
  wire [64:0] _by_divide_num_T_1 = regs_0[127:63]; // @[hard_cal.scala 91:58]
  wire [64:0] _by_divide_num_T_4 = {1'h0,regs_1[63:0]}; // @[hard_cal.scala 91:103]
  wire [64:0] by_divide_num = $signed(_by_divide_num_T_1) - $signed(_by_divide_num_T_4); // @[hard_cal.scala 91:65]
  wire  minus_answer = $signed(by_divide_num) >= 65'sh0; // @[hard_cal.scala 92:35]
  wire [64:0] _regs0_to_be_T = $signed(_by_divide_num_T_1) - $signed(_by_divide_num_T_4); // @[hard_cal.scala 93:58]
  wire [63:0] _regs0_to_be_T_3 = minus_answer ? _regs0_to_be_T[63:0] : regs_0[126:63]; // @[hard_cal.scala 93:30]
  wire [127:0] regs0_to_be = {_regs0_to_be_T_3,regs_0[62:0],1'h0}; // @[Cat.scala 31:58]
  wire [64:0] _result_reg_T = {result_reg, 1'h0}; // @[hard_cal.scala 97:49]
  wire [63:0] _result_reg_T_2 = {_result_reg_T[63:1],minus_answer}; // @[Cat.scala 31:58]
  wire [63:0] _io_result_0_T = ~_result_reg_T_2; // @[hard_cal.scala 103:38]
  wire [63:0] _io_result_0_T_2 = _io_result_0_T + 64'h1; // @[hard_cal.scala 103:60]
  wire [63:0] _io_result_1_T = ~_regs0_to_be_T_3; // @[hard_cal.scala 103:38]
  wire [63:0] _io_result_1_T_2 = _io_result_1_T + 64'h1; // @[hard_cal.scala 103:60]
  wire [6:0] _io_Output_valid_T_1 = 7'h40 - 7'h1; // @[hard_cal.scala 105:45]
  assign io_result_0 = result_sign_0 ? _io_result_0_T_2 : _result_reg_T_2; // @[hard_cal.scala 103:17]
  assign io_result_1 = result_sign_1 ? _io_result_1_T_2 : _regs0_to_be_T_3; // @[hard_cal.scala 103:17]
  assign io_input_ready = ~cal_start; // @[hard_cal.scala 106:23]
  assign io_Output_valid = counter == _io_Output_valid_T_1; // @[hard_cal.scala 105:33]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 94:19]
      regs_0 <= 128'h0;
    end else if (_cal_start_T) begin // @[hard_cal.scala 94:67]
      regs_0 <= {{64'd0}, data_in_0};
    end else if (cal_start) begin
      regs_0 <= regs0_to_be;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 96:19]
      regs_1 <= 128'h0;
    end else if (_cal_start_T) begin
      regs_1 <= {{64'd0}, data_in_1};
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 68:19]
      counter <= 7'h0;
    end else if (cal_start) begin
      counter <= _counter_T_1;
    end else begin
      counter <= 7'h0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 67:21]
      cal_start <= 1'h0;
    end else begin
      cal_start <= io_input_valid & io_input_ready | _cal_start_T_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 97:22]
      result_reg <= 64'h0;
    end else if (cal_start) begin
      result_reg <= _result_reg_T_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  regs_0 = _RAND_0[127:0];
  _RAND_1 = {4{`RANDOM}};
  regs_1 = _RAND_1[127:0];
  _RAND_2 = {1{`RANDOM}};
  counter = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  cal_start = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  result_reg = _RAND_4[63:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    regs_0 = 128'h0;
  end
  if (reset) begin
    regs_1 = 128'h0;
  end
  if (reset) begin
    counter = 7'h0;
  end
  if (reset) begin
    cal_start = 1'h0;
  end
  if (reset) begin
    result_reg = 64'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module div_simple_1(
  input         clock,
  input         reset,
  output [31:0] io_result_0,
  output [31:0] io_result_1,
  input  [31:0] io_data_0,
  input  [31:0] io_data_1,
  input         io_input_valid,
  output        io_input_ready,
  output        io_Output_valid,
  input         io_signed
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] regs_0; // @[hard_cal.scala 63:23]
  reg [63:0] regs_1; // @[hard_cal.scala 63:23]
  reg [5:0] counter; // @[hard_cal.scala 65:26]
  reg  cal_start; // @[hard_cal.scala 66:28]
  wire  _cal_start_T = io_input_valid & io_input_ready; // @[hard_cal.scala 67:37]
  wire  _cal_start_T_2 = counter == 6'h20 ? 1'h0 : cal_start; // @[hard_cal.scala 67:69]
  wire [5:0] _counter_T_1 = counter + 6'h1; // @[hard_cal.scala 68:39]
  reg [31:0] result_reg; // @[hard_cal.scala 70:29]
  wire [31:0] _data_in_0_T_2 = ~io_data_0; // @[hard_cal.scala 74:59]
  wire [31:0] _data_in_0_T_4 = _data_in_0_T_2 + 32'h1; // @[hard_cal.scala 74:76]
  wire [31:0] data_in_0 = io_signed & io_data_0[31] ? _data_in_0_T_4 : io_data_0; // @[hard_cal.scala 74:17]
  wire [31:0] _data_in_1_T_2 = ~io_data_1; // @[hard_cal.scala 74:59]
  wire [31:0] _data_in_1_T_4 = _data_in_1_T_2 + 32'h1; // @[hard_cal.scala 74:76]
  wire [31:0] data_in_1 = io_signed & io_data_1[31] ? _data_in_1_T_4 : io_data_1; // @[hard_cal.scala 74:17]
  wire [1:0] _T_2 = {io_data_0[31],io_data_1[31]}; // @[Cat.scala 31:58]
  wire  _T_6_1 = 2'h1 == _T_2 ? 1'h0 : 1'h1; // @[Mux.scala 81:58]
  wire  _T_8_0 = 2'h0 == _T_2 ? 1'h0 : 2'h1 == _T_2 | 2'h2 == _T_2; // @[Mux.scala 81:58]
  wire  _T_8_1 = 2'h0 == _T_2 ? 1'h0 : _T_6_1; // @[Mux.scala 81:58]
  wire  result_sign_0 = io_signed & _T_8_0; // @[hard_cal.scala 77:23]
  wire  result_sign_1 = io_signed & _T_8_1; // @[hard_cal.scala 77:23]
  wire [32:0] _by_divide_num_T_1 = regs_0[63:31]; // @[hard_cal.scala 91:58]
  wire [32:0] _by_divide_num_T_4 = {1'h0,regs_1[31:0]}; // @[hard_cal.scala 91:103]
  wire [32:0] by_divide_num = $signed(_by_divide_num_T_1) - $signed(_by_divide_num_T_4); // @[hard_cal.scala 91:65]
  wire  minus_answer = $signed(by_divide_num) >= 33'sh0; // @[hard_cal.scala 92:35]
  wire [32:0] _regs0_to_be_T = $signed(_by_divide_num_T_1) - $signed(_by_divide_num_T_4); // @[hard_cal.scala 93:58]
  wire [31:0] _regs0_to_be_T_3 = minus_answer ? _regs0_to_be_T[31:0] : regs_0[62:31]; // @[hard_cal.scala 93:30]
  wire [63:0] regs0_to_be = {_regs0_to_be_T_3,regs_0[30:0],1'h0}; // @[Cat.scala 31:58]
  wire [32:0] _result_reg_T = {result_reg, 1'h0}; // @[hard_cal.scala 97:49]
  wire [31:0] _result_reg_T_2 = {_result_reg_T[31:1],minus_answer}; // @[Cat.scala 31:58]
  wire [31:0] _io_result_0_T = ~_result_reg_T_2; // @[hard_cal.scala 103:38]
  wire [31:0] _io_result_0_T_2 = _io_result_0_T + 32'h1; // @[hard_cal.scala 103:60]
  wire [31:0] _io_result_1_T = ~_regs0_to_be_T_3; // @[hard_cal.scala 103:38]
  wire [31:0] _io_result_1_T_2 = _io_result_1_T + 32'h1; // @[hard_cal.scala 103:60]
  wire [5:0] _io_Output_valid_T_1 = 6'h20 - 6'h1; // @[hard_cal.scala 105:45]
  assign io_result_0 = result_sign_0 ? _io_result_0_T_2 : _result_reg_T_2; // @[hard_cal.scala 103:17]
  assign io_result_1 = result_sign_1 ? _io_result_1_T_2 : _regs0_to_be_T_3; // @[hard_cal.scala 103:17]
  assign io_input_ready = ~cal_start; // @[hard_cal.scala 106:23]
  assign io_Output_valid = counter == _io_Output_valid_T_1; // @[hard_cal.scala 105:33]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 94:19]
      regs_0 <= 64'h0;
    end else if (_cal_start_T) begin // @[hard_cal.scala 94:67]
      regs_0 <= {{32'd0}, data_in_0};
    end else if (cal_start) begin
      regs_0 <= regs0_to_be;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 96:19]
      regs_1 <= 64'h0;
    end else if (_cal_start_T) begin
      regs_1 <= {{32'd0}, data_in_1};
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 68:19]
      counter <= 6'h0;
    end else if (cal_start) begin
      counter <= _counter_T_1;
    end else begin
      counter <= 6'h0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 67:21]
      cal_start <= 1'h0;
    end else begin
      cal_start <= io_input_valid & io_input_ready | _cal_start_T_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[hard_cal.scala 97:22]
      result_reg <= 32'h0;
    end else if (cal_start) begin
      result_reg <= _result_reg_T_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  regs_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  regs_1 = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  counter = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  cal_start = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  result_reg = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    regs_0 = 64'h0;
  end
  if (reset) begin
    regs_1 = 64'h0;
  end
  if (reset) begin
    counter = 6'h0;
  end
  if (reset) begin
    cal_start = 1'h0;
  end
  if (reset) begin
    result_reg = 32'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module muldiv(
  input         clock,
  input         reset,
  input         io_en,
  input  [23:0] io_ctrl,
  input  [63:0] io_in1,
  input  [63:0] io_in2,
  output [63:0] io_data_out,
  output        io_pending
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  mul_hard_clock; // @[muldiv.scala 356:32]
  wire  mul_hard_reset; // @[muldiv.scala 356:32]
  wire [65:0] mul_hard_io_result_0; // @[muldiv.scala 356:32]
  wire [65:0] mul_hard_io_result_1; // @[muldiv.scala 356:32]
  wire [65:0] mul_hard_io_data_0; // @[muldiv.scala 356:32]
  wire [65:0] mul_hard_io_data_1; // @[muldiv.scala 356:32]
  wire  mul_hard_io_input_valid; // @[muldiv.scala 356:32]
  wire  mul_hard_io_input_ready; // @[muldiv.scala 356:32]
  wire  mul_hard_io_Output_valid; // @[muldiv.scala 356:32]
  wire  mul_hard_1_clock; // @[muldiv.scala 357:39]
  wire  mul_hard_1_reset; // @[muldiv.scala 357:39]
  wire [33:0] mul_hard_1_io_result_0; // @[muldiv.scala 357:39]
  wire [33:0] mul_hard_1_io_data_0; // @[muldiv.scala 357:39]
  wire [33:0] mul_hard_1_io_data_1; // @[muldiv.scala 357:39]
  wire  mul_hard_1_io_input_valid; // @[muldiv.scala 357:39]
  wire  mul_hard_1_io_input_ready; // @[muldiv.scala 357:39]
  wire  mul_hard_1_io_Output_valid; // @[muldiv.scala 357:39]
  wire  div_simple_clock; // @[muldiv.scala 385:32]
  wire  div_simple_reset; // @[muldiv.scala 385:32]
  wire [63:0] div_simple_io_result_0; // @[muldiv.scala 385:32]
  wire [63:0] div_simple_io_result_1; // @[muldiv.scala 385:32]
  wire [63:0] div_simple_io_data_0; // @[muldiv.scala 385:32]
  wire [63:0] div_simple_io_data_1; // @[muldiv.scala 385:32]
  wire  div_simple_io_input_valid; // @[muldiv.scala 385:32]
  wire  div_simple_io_input_ready; // @[muldiv.scala 385:32]
  wire  div_simple_io_Output_valid; // @[muldiv.scala 385:32]
  wire  div_simple_io_signed; // @[muldiv.scala 385:32]
  wire  div_simple_1_clock; // @[muldiv.scala 386:39]
  wire  div_simple_1_reset; // @[muldiv.scala 386:39]
  wire [31:0] div_simple_1_io_result_0; // @[muldiv.scala 386:39]
  wire [31:0] div_simple_1_io_result_1; // @[muldiv.scala 386:39]
  wire [31:0] div_simple_1_io_data_0; // @[muldiv.scala 386:39]
  wire [31:0] div_simple_1_io_data_1; // @[muldiv.scala 386:39]
  wire  div_simple_1_io_input_valid; // @[muldiv.scala 386:39]
  wire  div_simple_1_io_input_ready; // @[muldiv.scala 386:39]
  wire  div_simple_1_io_Output_valid; // @[muldiv.scala 386:39]
  wire  div_simple_1_io_signed; // @[muldiv.scala 386:39]
  wire [23:0] _cal_mul_T_1 = {{9'd0}, io_ctrl[23:9]}; // @[muldiv.scala 300:48]
  wire [23:0] _cal_mul_T_3 = {{12'd0}, io_ctrl[23:12]}; // @[muldiv.scala 300:71]
  wire [23:0] _cal_mul_T_6 = {{10'd0}, io_ctrl[23:10]}; // @[muldiv.scala 301:20]
  wire  _cal_mul_T_8 = _cal_mul_T_1[0] | _cal_mul_T_3[0] | _cal_mul_T_6[0]; // @[muldiv.scala 300:87]
  wire [23:0] _cal_mul_T_9 = {{11'd0}, io_ctrl[23:11]}; // @[muldiv.scala 301:46]
  wire  _cal_mul_T_11 = _cal_mul_T_8 | _cal_mul_T_9[0]; // @[muldiv.scala 301:36]
  wire  cal_mul = io_en & _cal_mul_T_11; // @[muldiv.scala 300:34]
  wire [23:0] _cal_div_T_1 = {{1'd0}, io_ctrl[23:1]}; // @[muldiv.scala 302:48]
  wire [23:0] _cal_div_T_6 = {{3'd0}, io_ctrl[23:3]}; // @[muldiv.scala 303:21]
  wire  _cal_div_T_8 = _cal_div_T_1[0] | io_ctrl[0] | _cal_div_T_6[0]; // @[muldiv.scala 302:85]
  wire [23:0] _cal_div_T_9 = {{2'd0}, io_ctrl[23:2]}; // @[muldiv.scala 303:45]
  wire  _cal_div_T_11 = _cal_div_T_8 | _cal_div_T_9[0]; // @[muldiv.scala 303:35]
  wire  cal_div = io_en & _cal_div_T_11; // @[muldiv.scala 302:34]
  wire [23:0] _cal_divw_T_1 = {{4'd0}, io_ctrl[23:4]}; // @[muldiv.scala 304:44]
  wire [23:0] _cal_divw_T_3 = {{5'd0}, io_ctrl[23:5]}; // @[muldiv.scala 304:69]
  wire [23:0] _cal_divw_T_6 = {{6'd0}, io_ctrl[23:6]}; // @[muldiv.scala 304:99]
  wire [23:0] _cal_divw_T_9 = {{7'd0}, io_ctrl[23:7]}; // @[muldiv.scala 304:125]
  wire  cal_divw = io_en & (_cal_divw_T_1[0] | _cal_divw_T_3[0] | _cal_divw_T_6[0] | _cal_divw_T_9[0]); // @[muldiv.scala 304:33]
  wire [23:0] _cal_mulw_T_1 = {{8'd0}, io_ctrl[23:8]}; // @[muldiv.scala 305:45]
  wire  cal_mulw = io_en & _cal_mulw_T_1[0]; // @[muldiv.scala 305:33]
  reg [3:0] work_state; // @[muldiv.scala 308:30]
  reg [23:0] ctrl_data; // @[muldiv.scala 315:28]
  wire  _work_state_T = work_state == 4'h0; // @[muldiv.scala 317:34]
  wire  _work_state_T_1 = cal_mul & work_state == 4'h0; // @[muldiv.scala 317:20]
  wire  _work_state_T_3 = cal_mulw & _work_state_T; // @[muldiv.scala 318:20]
  wire  _work_state_T_5 = cal_div & _work_state_T; // @[muldiv.scala 319:20]
  wire  _work_state_T_7 = cal_divw & _work_state_T; // @[muldiv.scala 320:20]
  wire  _work_state_T_8 = work_state == 4'h1; // @[muldiv.scala 321:37]
  wire  _work_state_T_9 = work_state == 4'h2; // @[muldiv.scala 321:69]
  wire  _cal_end_mul_T_1 = _work_state_T_8 & mul_hard_io_Output_valid; // @[muldiv.scala 368:43]
  wire  _cal_end_mul_T_3 = _work_state_T_9 & mul_hard_1_io_Output_valid; // @[muldiv.scala 369:44]
  wire  cal_end_mul = _cal_end_mul_T_1 | _cal_end_mul_T_3; // @[Mux.scala 101:16]
  wire  _work_state_T_11 = cal_end_mul & (work_state == 4'h1 | work_state == 4'h2); // @[muldiv.scala 321:22]
  wire  _work_state_T_12 = work_state == 4'h3; // @[muldiv.scala 322:38]
  wire  _work_state_T_13 = work_state == 4'h5; // @[muldiv.scala 322:70]
  wire  _cal_end_div_T_1 = _work_state_T_12 & div_simple_io_Output_valid; // @[muldiv.scala 397:43]
  wire  _cal_end_div_T_3 = _work_state_T_13 & div_simple_1_io_Output_valid; // @[muldiv.scala 398:44]
  wire  cal_end_div = _cal_end_div_T_1 | _cal_end_div_T_3; // @[Mux.scala 101:16]
  wire  _work_state_T_15 = cal_end_div & (work_state == 4'h3 | work_state == 4'h5); // @[muldiv.scala 322:23]
  wire  _work_state_T_16 = work_state == 4'h4; // @[muldiv.scala 323:21]
  wire [3:0] _work_state_T_17 = _work_state_T_16 ? 4'h0 : work_state; // @[Mux.scala 101:16]
  wire [3:0] _work_state_T_18 = _work_state_T_15 ? 4'h4 : _work_state_T_17; // @[Mux.scala 101:16]
  wire [3:0] _work_state_T_19 = _work_state_T_11 ? 4'h4 : _work_state_T_18; // @[Mux.scala 101:16]
  wire  cal_signed = _cal_mul_T_1[0] | _cal_mul_T_6[0] | _cal_mulw_T_1[0] | _cal_mul_T_3[0]; // @[muldiv.scala 358:95]
  wire [65:0] _T_4 = {io_in1[63],io_in1[63],io_in1}; // @[Cat.scala 31:58]
  wire [64:0] _T_6 = {1'h0,io_in1}; // @[Cat.scala 31:58]
  wire [65:0] _T_12 = {io_in2[63],io_in2[63],io_in2}; // @[Cat.scala 31:58]
  wire [64:0] _T_14 = {1'h0,io_in2}; // @[Cat.scala 31:58]
  wire [33:0] _T_21 = {io_in1[31],io_in1[31],io_in1[31:0]}; // @[Cat.scala 31:58]
  wire [32:0] _T_24 = {1'h0,io_in1[31:0]}; // @[Cat.scala 31:58]
  wire [33:0] _T_31 = {io_in2[31],io_in2[31],io_in2[31:0]}; // @[Cat.scala 31:58]
  wire [32:0] _T_34 = {1'h0,io_in2[31:0]}; // @[Cat.scala 31:58]
  wire [131:0] final_result = {mul_hard_io_result_1,mul_hard_io_result_0}; // @[Cat.scala 31:58]
  reg [63:0] mul_cal_reg; // @[muldiv.scala 372:34]
  wire [23:0] _access_mul_result_T = {{9'd0}, ctrl_data[23:9]}; // @[muldiv.scala 374:30]
  wire [23:0] _access_mul_result_T_3 = {{10'd0}, ctrl_data[23:10]}; // @[muldiv.scala 375:30]
  wire [23:0] _access_mul_result_T_6 = {{11'd0}, ctrl_data[23:11]}; // @[muldiv.scala 376:30]
  wire [23:0] _access_mul_result_T_9 = {{12'd0}, ctrl_data[23:12]}; // @[muldiv.scala 377:30]
  wire [23:0] _access_mul_result_T_12 = {{8'd0}, ctrl_data[23:8]}; // @[muldiv.scala 378:30]
  wire [7:0] access_mul_result_lo_lo = {mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31]
    ,mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],
    mul_hard_1_io_result_0[31]}; // @[Cat.scala 31:58]
  wire [15:0] access_mul_result_lo = {mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],
    mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],
    mul_hard_1_io_result_0[31],access_mul_result_lo_lo}; // @[Cat.scala 31:58]
  wire [31:0] _access_mul_result_T_47 = {mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31
    ],mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],mul_hard_1_io_result_0[31],
    mul_hard_1_io_result_0[31],access_mul_result_lo_lo,access_mul_result_lo}; // @[Cat.scala 31:58]
  wire [63:0] _access_mul_result_T_49 = {_access_mul_result_T_47,mul_hard_1_io_result_0[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _access_mul_result_T_50 = _access_mul_result_T[0] ? final_result[63:0] : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_mul_result_T_51 = _access_mul_result_T_3[0] ? final_result[127:64] : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_mul_result_T_52 = _access_mul_result_T_6[0] ? final_result[127:64] : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_mul_result_T_53 = _access_mul_result_T_9[0] ? final_result[127:64] : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_mul_result_T_54 = _access_mul_result_T_12[0] ? _access_mul_result_T_49 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_mul_result_T_55 = _access_mul_result_T_50 | _access_mul_result_T_51; // @[Mux.scala 27:73]
  wire [63:0] _access_mul_result_T_56 = _access_mul_result_T_55 | _access_mul_result_T_52; // @[Mux.scala 27:73]
  wire [63:0] _access_mul_result_T_57 = _access_mul_result_T_56 | _access_mul_result_T_53; // @[Mux.scala 27:73]
  wire [63:0] access_mul_result = _access_mul_result_T_57 | _access_mul_result_T_54; // @[Mux.scala 27:73]
  wire [63:0] cal_mul_result = cal_end_mul ? access_mul_result : mul_cal_reg; // @[muldiv.scala 380:30]
  reg [63:0] div_cal_reg; // @[muldiv.scala 400:34]
  wire [23:0] _access_div_result_T = {{1'd0}, ctrl_data[23:1]}; // @[muldiv.scala 402:30]
  wire [23:0] _access_div_result_T_4 = {{3'd0}, ctrl_data[23:3]}; // @[muldiv.scala 404:30]
  wire [23:0] _access_div_result_T_6 = {{2'd0}, ctrl_data[23:2]}; // @[muldiv.scala 405:30]
  wire [23:0] _access_div_result_T_8 = {{4'd0}, ctrl_data[23:4]}; // @[muldiv.scala 406:30]
  wire [7:0] access_div_result_lo_lo = {div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],
    div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],
    div_simple_1_io_result_0[31],div_simple_1_io_result_0[31]}; // @[Cat.scala 31:58]
  wire [15:0] access_div_result_lo = {div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],div_simple_1_io_result_0
    [31],div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],div_simple_1_io_result_0
    [31],div_simple_1_io_result_0[31],access_div_result_lo_lo}; // @[Cat.scala 31:58]
  wire [31:0] _access_div_result_T_42 = {div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],
    div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],
    div_simple_1_io_result_0[31],div_simple_1_io_result_0[31],access_div_result_lo_lo,access_div_result_lo}; // @[Cat.scala 31:58]
  wire [31:0] _access_div_result_T_43 = div_simple_1_io_result_0; // @[macros.scala 432:65]
  wire [63:0] _access_div_result_T_44 = {_access_div_result_T_42,_access_div_result_T_43}; // @[Cat.scala 31:58]
  wire [23:0] _access_div_result_T_45 = {{5'd0}, ctrl_data[23:5]}; // @[muldiv.scala 407:30]
  wire [23:0] _access_div_result_T_82 = {{6'd0}, ctrl_data[23:6]}; // @[muldiv.scala 408:30]
  wire [7:0] access_div_result_lo_lo_2 = {div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],
    div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],
    div_simple_1_io_result_1[31],div_simple_1_io_result_1[31]}; // @[Cat.scala 31:58]
  wire [15:0] access_div_result_lo_2 = {div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],
    div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],
    div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],access_div_result_lo_lo_2}; // @[Cat.scala 31:58]
  wire [31:0] _access_div_result_T_116 = {div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],
    div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],
    div_simple_1_io_result_1[31],div_simple_1_io_result_1[31],access_div_result_lo_lo_2,access_div_result_lo_2}; // @[Cat.scala 31:58]
  wire [31:0] _access_div_result_T_117 = div_simple_1_io_result_1; // @[macros.scala 432:65]
  wire [63:0] _access_div_result_T_118 = {_access_div_result_T_116,_access_div_result_T_117}; // @[Cat.scala 31:58]
  wire [23:0] _access_div_result_T_119 = {{7'd0}, ctrl_data[23:7]}; // @[muldiv.scala 409:30]
  wire [63:0] _access_div_result_T_156 = _access_div_result_T[0] ? div_simple_io_result_0 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_157 = ctrl_data[0] ? div_simple_io_result_0 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_158 = _access_div_result_T_4[0] ? div_simple_io_result_1 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_159 = _access_div_result_T_6[0] ? div_simple_io_result_1 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_160 = _access_div_result_T_8[0] ? _access_div_result_T_44 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_161 = _access_div_result_T_45[0] ? _access_div_result_T_44 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_162 = _access_div_result_T_82[0] ? _access_div_result_T_118 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_163 = _access_div_result_T_119[0] ? _access_div_result_T_118 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_164 = _access_div_result_T_156 | _access_div_result_T_157; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_165 = _access_div_result_T_164 | _access_div_result_T_158; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_166 = _access_div_result_T_165 | _access_div_result_T_159; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_167 = _access_div_result_T_166 | _access_div_result_T_160; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_168 = _access_div_result_T_167 | _access_div_result_T_161; // @[Mux.scala 27:73]
  wire [63:0] _access_div_result_T_169 = _access_div_result_T_168 | _access_div_result_T_162; // @[Mux.scala 27:73]
  wire [63:0] access_div_result = _access_div_result_T_169 | _access_div_result_T_163; // @[Mux.scala 27:73]
  wire [63:0] cal_div_result = cal_end_div ? access_div_result : div_cal_reg; // @[muldiv.scala 411:30]
  wire [63:0] _io_data_out_T_26 = _cal_div_T_1[0] ? cal_div_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_27 = io_ctrl[0] ? cal_div_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_28 = _cal_divw_T_1[0] ? cal_div_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_29 = _cal_divw_T_3[0] ? cal_div_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_30 = _cal_div_T_6[0] ? cal_div_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_31 = _cal_div_T_9[0] ? cal_div_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_32 = _cal_divw_T_6[0] ? cal_div_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_33 = _cal_divw_T_9[0] ? cal_div_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_34 = _cal_mul_T_1[0] ? cal_mul_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_35 = _cal_mulw_T_1[0] ? cal_mul_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_36 = _cal_mul_T_6[0] ? cal_mul_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_37 = _cal_mul_T_9[0] ? cal_mul_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_38 = _cal_mul_T_3[0] ? cal_mul_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_39 = _io_data_out_T_26 | _io_data_out_T_27; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_40 = _io_data_out_T_39 | _io_data_out_T_28; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_41 = _io_data_out_T_40 | _io_data_out_T_29; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_42 = _io_data_out_T_41 | _io_data_out_T_30; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_43 = _io_data_out_T_42 | _io_data_out_T_31; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_44 = _io_data_out_T_43 | _io_data_out_T_32; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_45 = _io_data_out_T_44 | _io_data_out_T_33; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_46 = _io_data_out_T_45 | _io_data_out_T_34; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_47 = _io_data_out_T_46 | _io_data_out_T_35; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_48 = _io_data_out_T_47 | _io_data_out_T_36; // @[Mux.scala 27:73]
  wire [63:0] _io_data_out_T_49 = _io_data_out_T_48 | _io_data_out_T_37; // @[Mux.scala 27:73]
  mul_hard mul_hard ( // @[muldiv.scala 356:32]
    .clock(mul_hard_clock),
    .reset(mul_hard_reset),
    .io_result_0(mul_hard_io_result_0),
    .io_result_1(mul_hard_io_result_1),
    .io_data_0(mul_hard_io_data_0),
    .io_data_1(mul_hard_io_data_1),
    .io_input_valid(mul_hard_io_input_valid),
    .io_input_ready(mul_hard_io_input_ready),
    .io_Output_valid(mul_hard_io_Output_valid)
  );
  mul_hard_1 mul_hard_1 ( // @[muldiv.scala 357:39]
    .clock(mul_hard_1_clock),
    .reset(mul_hard_1_reset),
    .io_result_0(mul_hard_1_io_result_0),
    .io_data_0(mul_hard_1_io_data_0),
    .io_data_1(mul_hard_1_io_data_1),
    .io_input_valid(mul_hard_1_io_input_valid),
    .io_input_ready(mul_hard_1_io_input_ready),
    .io_Output_valid(mul_hard_1_io_Output_valid)
  );
  div_simple div_simple ( // @[muldiv.scala 385:32]
    .clock(div_simple_clock),
    .reset(div_simple_reset),
    .io_result_0(div_simple_io_result_0),
    .io_result_1(div_simple_io_result_1),
    .io_data_0(div_simple_io_data_0),
    .io_data_1(div_simple_io_data_1),
    .io_input_valid(div_simple_io_input_valid),
    .io_input_ready(div_simple_io_input_ready),
    .io_Output_valid(div_simple_io_Output_valid),
    .io_signed(div_simple_io_signed)
  );
  div_simple_1 div_simple_1 ( // @[muldiv.scala 386:39]
    .clock(div_simple_1_clock),
    .reset(div_simple_1_reset),
    .io_result_0(div_simple_1_io_result_0),
    .io_result_1(div_simple_1_io_result_1),
    .io_data_0(div_simple_1_io_data_0),
    .io_data_1(div_simple_1_io_data_1),
    .io_input_valid(div_simple_1_io_input_valid),
    .io_input_ready(div_simple_1_io_input_ready),
    .io_Output_valid(div_simple_1_io_Output_valid),
    .io_signed(div_simple_1_io_signed)
  );
  assign io_data_out = _io_data_out_T_49 | _io_data_out_T_38; // @[Mux.scala 27:73]
  assign io_pending = work_state != 4'h0 & work_state != 4'h4 | _work_state_T & (cal_mul | cal_mulw | cal_div | cal_divw
    ); // @[muldiv.scala 455:79]
  assign mul_hard_clock = clock;
  assign mul_hard_reset = reset;
  assign mul_hard_io_data_0 = cal_signed ? _T_4 : {{1'd0}, _T_6}; // @[muldiv.scala 361:34]
  assign mul_hard_io_data_1 = cal_signed ? _T_12 : {{1'd0}, _T_14}; // @[muldiv.scala 362:34]
  assign mul_hard_io_input_valid = _work_state_T & cal_mul; // @[muldiv.scala 365:66]
  assign mul_hard_1_clock = clock;
  assign mul_hard_1_reset = reset;
  assign mul_hard_1_io_data_0 = cal_signed ? _T_21 : {{1'd0}, _T_24}; // @[muldiv.scala 363:41]
  assign mul_hard_1_io_data_1 = cal_signed ? _T_31 : {{1'd0}, _T_34}; // @[muldiv.scala 364:41]
  assign mul_hard_1_io_input_valid = _work_state_T & cal_mulw; // @[muldiv.scala 366:72]
  assign div_simple_clock = clock;
  assign div_simple_reset = reset;
  assign div_simple_io_data_0 = io_in1; // @[muldiv.scala 390:28]
  assign div_simple_io_data_1 = io_in2; // @[muldiv.scala 391:28]
  assign div_simple_io_input_valid = _work_state_T & cal_div; // @[muldiv.scala 394:66]
  assign div_simple_io_signed = _cal_div_T_1[0] | _cal_divw_T_1[0] | _cal_div_T_6[0] | _cal_divw_T_6[0]; // @[muldiv.scala 387:96]
  assign div_simple_1_clock = clock;
  assign div_simple_1_reset = reset;
  assign div_simple_1_io_data_0 = io_in1[31:0]; // @[muldiv.scala 392:35]
  assign div_simple_1_io_data_1 = io_in2[31:0]; // @[muldiv.scala 393:35]
  assign div_simple_1_io_input_valid = _work_state_T & cal_divw; // @[muldiv.scala 395:72]
  assign div_simple_1_io_signed = _cal_div_T_1[0] | _cal_divw_T_1[0] | _cal_div_T_6[0] | _cal_divw_T_6[0]; // @[muldiv.scala 387:96]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Mux.scala 101:16]
      work_state <= 4'h0;
    end else if (_work_state_T_1) begin // @[Mux.scala 101:16]
      work_state <= 4'h1;
    end else if (_work_state_T_3) begin // @[Mux.scala 101:16]
      work_state <= 4'h2;
    end else if (_work_state_T_5) begin // @[Mux.scala 101:16]
      work_state <= 4'h3;
    end else if (_work_state_T_7) begin
      work_state <= 4'h5;
    end else begin
      work_state <= _work_state_T_19;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[muldiv.scala 325:22]
      ctrl_data <= 24'h0;
    end else if (_work_state_T) begin
      ctrl_data <= io_ctrl;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[muldiv.scala 381:27]
      mul_cal_reg <= 64'h0;
    end else if (cal_end_mul) begin
      mul_cal_reg <= access_mul_result;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[muldiv.scala 412:27]
      div_cal_reg <= 64'h0;
    end else if (cal_end_div) begin
      div_cal_reg <= access_div_result;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  work_state = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  ctrl_data = _RAND_1[23:0];
  _RAND_2 = {2{`RANDOM}};
  mul_cal_reg = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  div_cal_reg = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    work_state = 4'h0;
  end
  if (reset) begin
    ctrl_data = 24'h0;
  end
  if (reset) begin
    mul_cal_reg = 64'h0;
  end
  if (reset) begin
    div_cal_reg = 64'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module regfile(
  input           clock,
  input           reset,
  input  [4:0]    io_A1,
  input  [4:0]    io_A2,
  input           io_WE3,
  input  [4:0]    io_A3,
  input  [63:0]   io_WD3,
  output [63:0]   io_RD1,
  output [63:0]   io_RD2,
  output [2047:0] io_reg_file_alL_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] regs_0; // @[regfile.scala 24:23]
  reg [63:0] regs_1; // @[regfile.scala 24:23]
  reg [63:0] regs_2; // @[regfile.scala 24:23]
  reg [63:0] regs_3; // @[regfile.scala 24:23]
  reg [63:0] regs_4; // @[regfile.scala 24:23]
  reg [63:0] regs_5; // @[regfile.scala 24:23]
  reg [63:0] regs_6; // @[regfile.scala 24:23]
  reg [63:0] regs_7; // @[regfile.scala 24:23]
  reg [63:0] regs_8; // @[regfile.scala 24:23]
  reg [63:0] regs_9; // @[regfile.scala 24:23]
  reg [63:0] regs_10; // @[regfile.scala 24:23]
  reg [63:0] regs_11; // @[regfile.scala 24:23]
  reg [63:0] regs_12; // @[regfile.scala 24:23]
  reg [63:0] regs_13; // @[regfile.scala 24:23]
  reg [63:0] regs_14; // @[regfile.scala 24:23]
  reg [63:0] regs_15; // @[regfile.scala 24:23]
  reg [63:0] regs_16; // @[regfile.scala 24:23]
  reg [63:0] regs_17; // @[regfile.scala 24:23]
  reg [63:0] regs_18; // @[regfile.scala 24:23]
  reg [63:0] regs_19; // @[regfile.scala 24:23]
  reg [63:0] regs_20; // @[regfile.scala 24:23]
  reg [63:0] regs_21; // @[regfile.scala 24:23]
  reg [63:0] regs_22; // @[regfile.scala 24:23]
  reg [63:0] regs_23; // @[regfile.scala 24:23]
  reg [63:0] regs_24; // @[regfile.scala 24:23]
  reg [63:0] regs_25; // @[regfile.scala 24:23]
  reg [63:0] regs_26; // @[regfile.scala 24:23]
  reg [63:0] regs_27; // @[regfile.scala 24:23]
  reg [63:0] regs_28; // @[regfile.scala 24:23]
  reg [63:0] regs_29; // @[regfile.scala 24:23]
  reg [63:0] regs_30; // @[regfile.scala 24:23]
  reg [63:0] regs_31; // @[regfile.scala 24:23]
  wire [63:0] _GEN_1 = 5'h1 == io_A3 ? regs_1 : regs_0; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_2 = 5'h2 == io_A3 ? regs_2 : _GEN_1; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_3 = 5'h3 == io_A3 ? regs_3 : _GEN_2; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_4 = 5'h4 == io_A3 ? regs_4 : _GEN_3; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_5 = 5'h5 == io_A3 ? regs_5 : _GEN_4; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_6 = 5'h6 == io_A3 ? regs_6 : _GEN_5; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_7 = 5'h7 == io_A3 ? regs_7 : _GEN_6; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_8 = 5'h8 == io_A3 ? regs_8 : _GEN_7; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_9 = 5'h9 == io_A3 ? regs_9 : _GEN_8; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_10 = 5'ha == io_A3 ? regs_10 : _GEN_9; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_11 = 5'hb == io_A3 ? regs_11 : _GEN_10; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_12 = 5'hc == io_A3 ? regs_12 : _GEN_11; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_13 = 5'hd == io_A3 ? regs_13 : _GEN_12; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_14 = 5'he == io_A3 ? regs_14 : _GEN_13; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_15 = 5'hf == io_A3 ? regs_15 : _GEN_14; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_16 = 5'h10 == io_A3 ? regs_16 : _GEN_15; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_17 = 5'h11 == io_A3 ? regs_17 : _GEN_16; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_18 = 5'h12 == io_A3 ? regs_18 : _GEN_17; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_19 = 5'h13 == io_A3 ? regs_19 : _GEN_18; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_20 = 5'h14 == io_A3 ? regs_20 : _GEN_19; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_21 = 5'h15 == io_A3 ? regs_21 : _GEN_20; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_22 = 5'h16 == io_A3 ? regs_22 : _GEN_21; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_23 = 5'h17 == io_A3 ? regs_23 : _GEN_22; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_24 = 5'h18 == io_A3 ? regs_24 : _GEN_23; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_25 = 5'h19 == io_A3 ? regs_25 : _GEN_24; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_26 = 5'h1a == io_A3 ? regs_26 : _GEN_25; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_27 = 5'h1b == io_A3 ? regs_27 : _GEN_26; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_28 = 5'h1c == io_A3 ? regs_28 : _GEN_27; // @[regfile.scala 26:{23,23}]
  wire [63:0] _GEN_29 = 5'h1d == io_A3 ? regs_29 : _GEN_28; // @[regfile.scala 26:{23,23}]
  wire [511:0] io_reg_file_alL_out_lo_lo = {regs_7,regs_6,regs_5,regs_4,regs_3,regs_2,regs_1,regs_0}; // @[Cat.scala 31:58]
  wire [1023:0] io_reg_file_alL_out_lo = {regs_15,regs_14,regs_13,regs_12,regs_11,regs_10,regs_9,regs_8,
    io_reg_file_alL_out_lo_lo}; // @[Cat.scala 31:58]
  wire [511:0] io_reg_file_alL_out_hi_lo = {regs_23,regs_22,regs_21,regs_20,regs_19,regs_18,regs_17,regs_16}; // @[Cat.scala 31:58]
  wire [1023:0] io_reg_file_alL_out_hi = {regs_31,regs_30,regs_29,regs_28,regs_27,regs_26,regs_25,regs_24,
    io_reg_file_alL_out_hi_lo}; // @[Cat.scala 31:58]
  wire [63:0] _GEN_65 = 5'h1 == io_A1 ? regs_1 : regs_0; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_66 = 5'h2 == io_A1 ? regs_2 : _GEN_65; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_67 = 5'h3 == io_A1 ? regs_3 : _GEN_66; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_68 = 5'h4 == io_A1 ? regs_4 : _GEN_67; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_69 = 5'h5 == io_A1 ? regs_5 : _GEN_68; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_70 = 5'h6 == io_A1 ? regs_6 : _GEN_69; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_71 = 5'h7 == io_A1 ? regs_7 : _GEN_70; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_72 = 5'h8 == io_A1 ? regs_8 : _GEN_71; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_73 = 5'h9 == io_A1 ? regs_9 : _GEN_72; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_74 = 5'ha == io_A1 ? regs_10 : _GEN_73; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_75 = 5'hb == io_A1 ? regs_11 : _GEN_74; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_76 = 5'hc == io_A1 ? regs_12 : _GEN_75; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_77 = 5'hd == io_A1 ? regs_13 : _GEN_76; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_78 = 5'he == io_A1 ? regs_14 : _GEN_77; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_79 = 5'hf == io_A1 ? regs_15 : _GEN_78; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_80 = 5'h10 == io_A1 ? regs_16 : _GEN_79; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_81 = 5'h11 == io_A1 ? regs_17 : _GEN_80; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_82 = 5'h12 == io_A1 ? regs_18 : _GEN_81; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_83 = 5'h13 == io_A1 ? regs_19 : _GEN_82; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_84 = 5'h14 == io_A1 ? regs_20 : _GEN_83; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_85 = 5'h15 == io_A1 ? regs_21 : _GEN_84; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_86 = 5'h16 == io_A1 ? regs_22 : _GEN_85; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_87 = 5'h17 == io_A1 ? regs_23 : _GEN_86; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_88 = 5'h18 == io_A1 ? regs_24 : _GEN_87; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_89 = 5'h19 == io_A1 ? regs_25 : _GEN_88; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_90 = 5'h1a == io_A1 ? regs_26 : _GEN_89; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_91 = 5'h1b == io_A1 ? regs_27 : _GEN_90; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_92 = 5'h1c == io_A1 ? regs_28 : _GEN_91; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_93 = 5'h1d == io_A1 ? regs_29 : _GEN_92; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_94 = 5'h1e == io_A1 ? regs_30 : _GEN_93; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_95 = 5'h1f == io_A1 ? regs_31 : _GEN_94; // @[regfile.scala 31:{19,19}]
  wire [63:0] _GEN_97 = 5'h1 == io_A2 ? regs_1 : regs_0; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_98 = 5'h2 == io_A2 ? regs_2 : _GEN_97; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_99 = 5'h3 == io_A2 ? regs_3 : _GEN_98; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_100 = 5'h4 == io_A2 ? regs_4 : _GEN_99; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_101 = 5'h5 == io_A2 ? regs_5 : _GEN_100; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_102 = 5'h6 == io_A2 ? regs_6 : _GEN_101; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_103 = 5'h7 == io_A2 ? regs_7 : _GEN_102; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_104 = 5'h8 == io_A2 ? regs_8 : _GEN_103; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_105 = 5'h9 == io_A2 ? regs_9 : _GEN_104; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_106 = 5'ha == io_A2 ? regs_10 : _GEN_105; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_107 = 5'hb == io_A2 ? regs_11 : _GEN_106; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_108 = 5'hc == io_A2 ? regs_12 : _GEN_107; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_109 = 5'hd == io_A2 ? regs_13 : _GEN_108; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_110 = 5'he == io_A2 ? regs_14 : _GEN_109; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_111 = 5'hf == io_A2 ? regs_15 : _GEN_110; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_112 = 5'h10 == io_A2 ? regs_16 : _GEN_111; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_113 = 5'h11 == io_A2 ? regs_17 : _GEN_112; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_114 = 5'h12 == io_A2 ? regs_18 : _GEN_113; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_115 = 5'h13 == io_A2 ? regs_19 : _GEN_114; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_116 = 5'h14 == io_A2 ? regs_20 : _GEN_115; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_117 = 5'h15 == io_A2 ? regs_21 : _GEN_116; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_118 = 5'h16 == io_A2 ? regs_22 : _GEN_117; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_119 = 5'h17 == io_A2 ? regs_23 : _GEN_118; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_120 = 5'h18 == io_A2 ? regs_24 : _GEN_119; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_121 = 5'h19 == io_A2 ? regs_25 : _GEN_120; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_122 = 5'h1a == io_A2 ? regs_26 : _GEN_121; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_123 = 5'h1b == io_A2 ? regs_27 : _GEN_122; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_124 = 5'h1c == io_A2 ? regs_28 : _GEN_123; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_125 = 5'h1d == io_A2 ? regs_29 : _GEN_124; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_126 = 5'h1e == io_A2 ? regs_30 : _GEN_125; // @[regfile.scala 32:{19,19}]
  wire [63:0] _GEN_127 = 5'h1f == io_A2 ? regs_31 : _GEN_126; // @[regfile.scala 32:{19,19}]
  assign io_RD1 = io_WE3 & io_A1 == io_A3 & io_A1 != 5'h0 ? io_WD3 : _GEN_95; // @[regfile.scala 31:19]
  assign io_RD2 = io_WE3 & io_A2 == io_A3 & io_A2 != 5'h0 ? io_WD3 : _GEN_127; // @[regfile.scala 32:19]
  assign io_reg_file_alL_out = {io_reg_file_alL_out_hi,io_reg_file_alL_out_lo}; // @[Cat.scala 31:58]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_0 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h0 == io_A3) begin // @[regfile.scala 25:13]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_0 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_0 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_0 <= regs_30;
      end else begin
        regs_0 <= _GEN_29;
      end
    end else begin
      regs_0 <= 64'h0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_1 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h1 == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_1 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_1 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_1 <= regs_30;
      end else begin
        regs_1 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_2 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h2 == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_2 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_2 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_2 <= regs_30;
      end else begin
        regs_2 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_3 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h3 == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_3 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_3 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_3 <= regs_30;
      end else begin
        regs_3 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_4 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h4 == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_4 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_4 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_4 <= regs_30;
      end else begin
        regs_4 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_5 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h5 == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_5 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_5 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_5 <= regs_30;
      end else begin
        regs_5 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_6 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h6 == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_6 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_6 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_6 <= regs_30;
      end else begin
        regs_6 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_7 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h7 == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_7 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_7 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_7 <= regs_30;
      end else begin
        regs_7 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_8 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h8 == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_8 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_8 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_8 <= regs_30;
      end else begin
        regs_8 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_9 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h9 == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_9 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_9 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_9 <= regs_30;
      end else begin
        regs_9 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_10 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'ha == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_10 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_10 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_10 <= regs_30;
      end else begin
        regs_10 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_11 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'hb == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_11 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_11 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_11 <= regs_30;
      end else begin
        regs_11 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_12 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'hc == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_12 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_12 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_12 <= regs_30;
      end else begin
        regs_12 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_13 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'hd == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_13 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_13 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_13 <= regs_30;
      end else begin
        regs_13 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_14 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'he == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_14 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_14 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_14 <= regs_30;
      end else begin
        regs_14 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_15 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'hf == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_15 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_15 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_15 <= regs_30;
      end else begin
        regs_15 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_16 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h10 == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_16 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_16 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_16 <= regs_30;
      end else begin
        regs_16 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_17 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h11 == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_17 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_17 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_17 <= regs_30;
      end else begin
        regs_17 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_18 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h12 == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_18 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_18 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_18 <= regs_30;
      end else begin
        regs_18 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_19 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h13 == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_19 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_19 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_19 <= regs_30;
      end else begin
        regs_19 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_20 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h14 == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_20 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_20 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_20 <= regs_30;
      end else begin
        regs_20 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_21 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h15 == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_21 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_21 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_21 <= regs_30;
      end else begin
        regs_21 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_22 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h16 == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_22 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_22 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_22 <= regs_30;
      end else begin
        regs_22 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_23 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h17 == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_23 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_23 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_23 <= regs_30;
      end else begin
        regs_23 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_24 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h18 == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_24 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_24 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_24 <= regs_30;
      end else begin
        regs_24 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_25 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h19 == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_25 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_25 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_25 <= regs_30;
      end else begin
        regs_25 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_26 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h1a == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_26 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_26 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_26 <= regs_30;
      end else begin
        regs_26 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_27 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h1b == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_27 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_27 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_27 <= regs_30;
      end else begin
        regs_27 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_28 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h1c == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_28 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_28 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_28 <= regs_30;
      end else begin
        regs_28 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_29 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h1d == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_29 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_29 <= regs_31;
      end else if (5'h1e == io_A3) begin
        regs_29 <= regs_30;
      end else begin
        regs_29 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_30 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h1e == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_30 <= io_WD3;
      end else if (5'h1f == io_A3) begin
        regs_30 <= regs_31;
      end else if (!(5'h1e == io_A3)) begin
        regs_30 <= _GEN_29;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[regfile.scala 26:17]
      regs_31 <= 64'h0; // @[regfile.scala 26:{23,23,23,23,23}]
    end else if (5'h1f == io_A3) begin // @[regfile.scala 24:23]
      if (io_WE3 & io_A3 != 5'h0) begin
        regs_31 <= io_WD3;
      end else if (!(5'h1f == io_A3)) begin
        if (5'h1e == io_A3) begin
          regs_31 <= regs_30;
        end else begin
          regs_31 <= _GEN_29;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  regs_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  regs_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  regs_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  regs_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  regs_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  regs_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  regs_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  regs_7 = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  regs_8 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  regs_9 = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  regs_10 = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  regs_11 = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  regs_12 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  regs_13 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  regs_14 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  regs_15 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  regs_16 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  regs_17 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  regs_18 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  regs_19 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  regs_20 = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  regs_21 = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  regs_22 = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  regs_23 = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  regs_24 = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  regs_25 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  regs_26 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  regs_27 = _RAND_27[63:0];
  _RAND_28 = {2{`RANDOM}};
  regs_28 = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  regs_29 = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  regs_30 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  regs_31 = _RAND_31[63:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    regs_0 = 64'h0;
  end
  if (reset) begin
    regs_1 = 64'h0;
  end
  if (reset) begin
    regs_2 = 64'h0;
  end
  if (reset) begin
    regs_3 = 64'h0;
  end
  if (reset) begin
    regs_4 = 64'h0;
  end
  if (reset) begin
    regs_5 = 64'h0;
  end
  if (reset) begin
    regs_6 = 64'h0;
  end
  if (reset) begin
    regs_7 = 64'h0;
  end
  if (reset) begin
    regs_8 = 64'h0;
  end
  if (reset) begin
    regs_9 = 64'h0;
  end
  if (reset) begin
    regs_10 = 64'h0;
  end
  if (reset) begin
    regs_11 = 64'h0;
  end
  if (reset) begin
    regs_12 = 64'h0;
  end
  if (reset) begin
    regs_13 = 64'h0;
  end
  if (reset) begin
    regs_14 = 64'h0;
  end
  if (reset) begin
    regs_15 = 64'h0;
  end
  if (reset) begin
    regs_16 = 64'h0;
  end
  if (reset) begin
    regs_17 = 64'h0;
  end
  if (reset) begin
    regs_18 = 64'h0;
  end
  if (reset) begin
    regs_19 = 64'h0;
  end
  if (reset) begin
    regs_20 = 64'h0;
  end
  if (reset) begin
    regs_21 = 64'h0;
  end
  if (reset) begin
    regs_22 = 64'h0;
  end
  if (reset) begin
    regs_23 = 64'h0;
  end
  if (reset) begin
    regs_24 = 64'h0;
  end
  if (reset) begin
    regs_25 = 64'h0;
  end
  if (reset) begin
    regs_26 = 64'h0;
  end
  if (reset) begin
    regs_27 = 64'h0;
  end
  if (reset) begin
    regs_28 = 64'h0;
  end
  if (reset) begin
    regs_29 = 64'h0;
  end
  if (reset) begin
    regs_30 = 64'h0;
  end
  if (reset) begin
    regs_31 = 64'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Look_up_table_read_first_with_bundle(
  input         clock,
  input         reset,
  input  [3:0]  io_ar_addr,
  input  [3:0]  io_aw_addr,
  input         io_write,
  input  [63:0] io_in_pc,
  input  [31:0] io_in_inst,
  input  [63:0] io_in_pre_pc_target,
  input  [6:0]  io_in_pre_lookup_data,
  input  [3:0]  io_in_pre_hashcode,
  input  [1:0]  io_in_pre_pht,
  input  [6:0]  io_in_pre_bht,
  input  [7:0]  io_in_pre_lookup_value,
  input         io_in_pre_decoder_branchD_flag,
  input         io_in_pre_decoder_jump,
  input  [5:0]  io_in_pre_decoder_branchdata,
  input         io_in_pre_decoder_jr,
  input         io_in_true_branch_state,
  output [63:0] io_out_pc,
  output [31:0] io_out_inst,
  output [1:0]  io_out_exception_type,
  output [63:0] io_out_pre_pc_target,
  output [6:0]  io_out_pre_lookup_data,
  output [3:0]  io_out_pre_hashcode,
  output [1:0]  io_out_pre_pht,
  output [6:0]  io_out_pre_bht,
  output [7:0]  io_out_pre_lookup_value,
  output        io_out_pre_decoder_branchD_flag,
  output        io_out_pre_decoder_jump,
  output [5:0]  io_out_pre_decoder_branchdata,
  output        io_out_pre_decoder_jr,
  output        io_out_true_branch_state
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [63:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [63:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [63:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [63:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [63:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [63:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [63:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [63:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [63:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [63:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [63:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] btb_0_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_0_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_0_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_0_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_0_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_0_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_0_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_0_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg [7:0] btb_0_pre_lookup_value; // @[ports_lookup_table.scala 105:22]
  reg  btb_0_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_0_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_0_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_0_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_0_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_1_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_1_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_1_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_1_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_1_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_1_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_1_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_1_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg [7:0] btb_1_pre_lookup_value; // @[ports_lookup_table.scala 105:22]
  reg  btb_1_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_1_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_1_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_1_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_1_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_2_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_2_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_2_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_2_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_2_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_2_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_2_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_2_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg [7:0] btb_2_pre_lookup_value; // @[ports_lookup_table.scala 105:22]
  reg  btb_2_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_2_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_2_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_2_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_2_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_3_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_3_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_3_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_3_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_3_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_3_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_3_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_3_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg [7:0] btb_3_pre_lookup_value; // @[ports_lookup_table.scala 105:22]
  reg  btb_3_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_3_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_3_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_3_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_3_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_4_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_4_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_4_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_4_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_4_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_4_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_4_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_4_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg [7:0] btb_4_pre_lookup_value; // @[ports_lookup_table.scala 105:22]
  reg  btb_4_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_4_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_4_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_4_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_4_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_5_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_5_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_5_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_5_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_5_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_5_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_5_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_5_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg [7:0] btb_5_pre_lookup_value; // @[ports_lookup_table.scala 105:22]
  reg  btb_5_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_5_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_5_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_5_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_5_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_6_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_6_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_6_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_6_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_6_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_6_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_6_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_6_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg [7:0] btb_6_pre_lookup_value; // @[ports_lookup_table.scala 105:22]
  reg  btb_6_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_6_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_6_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_6_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_6_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_7_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_7_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_7_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_7_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_7_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_7_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_7_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_7_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg [7:0] btb_7_pre_lookup_value; // @[ports_lookup_table.scala 105:22]
  reg  btb_7_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_7_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_7_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_7_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_7_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_8_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_8_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_8_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_8_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_8_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_8_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_8_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_8_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg [7:0] btb_8_pre_lookup_value; // @[ports_lookup_table.scala 105:22]
  reg  btb_8_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_8_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_8_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_8_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_8_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_9_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_9_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_9_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_9_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_9_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_9_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_9_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_9_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg [7:0] btb_9_pre_lookup_value; // @[ports_lookup_table.scala 105:22]
  reg  btb_9_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_9_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_9_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_9_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_9_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_10_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_10_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_10_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_10_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_10_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_10_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_10_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_10_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg [7:0] btb_10_pre_lookup_value; // @[ports_lookup_table.scala 105:22]
  reg  btb_10_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_10_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_10_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_10_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_10_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_11_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_11_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_11_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_11_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_11_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_11_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_11_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_11_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg [7:0] btb_11_pre_lookup_value; // @[ports_lookup_table.scala 105:22]
  reg  btb_11_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_11_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_11_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_11_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_11_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_12_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_12_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_12_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_12_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_12_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_12_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_12_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_12_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg [7:0] btb_12_pre_lookup_value; // @[ports_lookup_table.scala 105:22]
  reg  btb_12_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_12_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_12_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_12_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_12_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_13_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_13_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_13_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_13_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_13_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_13_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_13_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_13_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg [7:0] btb_13_pre_lookup_value; // @[ports_lookup_table.scala 105:22]
  reg  btb_13_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_13_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_13_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_13_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_13_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_14_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_14_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_14_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_14_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_14_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_14_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_14_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_14_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg [7:0] btb_14_pre_lookup_value; // @[ports_lookup_table.scala 105:22]
  reg  btb_14_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_14_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_14_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_14_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_14_true_branch_state; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_15_pc; // @[ports_lookup_table.scala 105:22]
  reg [31:0] btb_15_inst; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_15_exception_type; // @[ports_lookup_table.scala 105:22]
  reg [63:0] btb_15_pre_pc_target; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_15_pre_lookup_data; // @[ports_lookup_table.scala 105:22]
  reg [3:0] btb_15_pre_hashcode; // @[ports_lookup_table.scala 105:22]
  reg [1:0] btb_15_pre_pht; // @[ports_lookup_table.scala 105:22]
  reg [6:0] btb_15_pre_bht; // @[ports_lookup_table.scala 105:22]
  reg [7:0] btb_15_pre_lookup_value; // @[ports_lookup_table.scala 105:22]
  reg  btb_15_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 105:22]
  reg  btb_15_pre_decoder_jump; // @[ports_lookup_table.scala 105:22]
  reg [5:0] btb_15_pre_decoder_branchdata; // @[ports_lookup_table.scala 105:22]
  reg  btb_15_pre_decoder_jr; // @[ports_lookup_table.scala 105:22]
  reg  btb_15_true_branch_state; // @[ports_lookup_table.scala 105:22]
  wire  _GEN_1 = 4'h1 == io_ar_addr ? btb_1_true_branch_state : btb_0_true_branch_state; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_2 = 4'h2 == io_ar_addr ? btb_2_true_branch_state : _GEN_1; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_3 = 4'h3 == io_ar_addr ? btb_3_true_branch_state : _GEN_2; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_4 = 4'h4 == io_ar_addr ? btb_4_true_branch_state : _GEN_3; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_5 = 4'h5 == io_ar_addr ? btb_5_true_branch_state : _GEN_4; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_6 = 4'h6 == io_ar_addr ? btb_6_true_branch_state : _GEN_5; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_7 = 4'h7 == io_ar_addr ? btb_7_true_branch_state : _GEN_6; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_8 = 4'h8 == io_ar_addr ? btb_8_true_branch_state : _GEN_7; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_9 = 4'h9 == io_ar_addr ? btb_9_true_branch_state : _GEN_8; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_10 = 4'ha == io_ar_addr ? btb_10_true_branch_state : _GEN_9; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_11 = 4'hb == io_ar_addr ? btb_11_true_branch_state : _GEN_10; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_12 = 4'hc == io_ar_addr ? btb_12_true_branch_state : _GEN_11; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_13 = 4'hd == io_ar_addr ? btb_13_true_branch_state : _GEN_12; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_14 = 4'he == io_ar_addr ? btb_14_true_branch_state : _GEN_13; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_17 = 4'h1 == io_ar_addr ? btb_1_pre_decoder_jr : btb_0_pre_decoder_jr; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_18 = 4'h2 == io_ar_addr ? btb_2_pre_decoder_jr : _GEN_17; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_19 = 4'h3 == io_ar_addr ? btb_3_pre_decoder_jr : _GEN_18; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_20 = 4'h4 == io_ar_addr ? btb_4_pre_decoder_jr : _GEN_19; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_21 = 4'h5 == io_ar_addr ? btb_5_pre_decoder_jr : _GEN_20; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_22 = 4'h6 == io_ar_addr ? btb_6_pre_decoder_jr : _GEN_21; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_23 = 4'h7 == io_ar_addr ? btb_7_pre_decoder_jr : _GEN_22; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_24 = 4'h8 == io_ar_addr ? btb_8_pre_decoder_jr : _GEN_23; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_25 = 4'h9 == io_ar_addr ? btb_9_pre_decoder_jr : _GEN_24; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_26 = 4'ha == io_ar_addr ? btb_10_pre_decoder_jr : _GEN_25; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_27 = 4'hb == io_ar_addr ? btb_11_pre_decoder_jr : _GEN_26; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_28 = 4'hc == io_ar_addr ? btb_12_pre_decoder_jr : _GEN_27; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_29 = 4'hd == io_ar_addr ? btb_13_pre_decoder_jr : _GEN_28; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_30 = 4'he == io_ar_addr ? btb_14_pre_decoder_jr : _GEN_29; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_33 = 4'h1 == io_ar_addr ? btb_1_pre_decoder_branchdata : btb_0_pre_decoder_branchdata; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_34 = 4'h2 == io_ar_addr ? btb_2_pre_decoder_branchdata : _GEN_33; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_35 = 4'h3 == io_ar_addr ? btb_3_pre_decoder_branchdata : _GEN_34; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_36 = 4'h4 == io_ar_addr ? btb_4_pre_decoder_branchdata : _GEN_35; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_37 = 4'h5 == io_ar_addr ? btb_5_pre_decoder_branchdata : _GEN_36; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_38 = 4'h6 == io_ar_addr ? btb_6_pre_decoder_branchdata : _GEN_37; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_39 = 4'h7 == io_ar_addr ? btb_7_pre_decoder_branchdata : _GEN_38; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_40 = 4'h8 == io_ar_addr ? btb_8_pre_decoder_branchdata : _GEN_39; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_41 = 4'h9 == io_ar_addr ? btb_9_pre_decoder_branchdata : _GEN_40; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_42 = 4'ha == io_ar_addr ? btb_10_pre_decoder_branchdata : _GEN_41; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_43 = 4'hb == io_ar_addr ? btb_11_pre_decoder_branchdata : _GEN_42; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_44 = 4'hc == io_ar_addr ? btb_12_pre_decoder_branchdata : _GEN_43; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_45 = 4'hd == io_ar_addr ? btb_13_pre_decoder_branchdata : _GEN_44; // @[ports_lookup_table.scala 106:{12,12}]
  wire [5:0] _GEN_46 = 4'he == io_ar_addr ? btb_14_pre_decoder_branchdata : _GEN_45; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_49 = 4'h1 == io_ar_addr ? btb_1_pre_decoder_jump : btb_0_pre_decoder_jump; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_50 = 4'h2 == io_ar_addr ? btb_2_pre_decoder_jump : _GEN_49; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_51 = 4'h3 == io_ar_addr ? btb_3_pre_decoder_jump : _GEN_50; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_52 = 4'h4 == io_ar_addr ? btb_4_pre_decoder_jump : _GEN_51; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_53 = 4'h5 == io_ar_addr ? btb_5_pre_decoder_jump : _GEN_52; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_54 = 4'h6 == io_ar_addr ? btb_6_pre_decoder_jump : _GEN_53; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_55 = 4'h7 == io_ar_addr ? btb_7_pre_decoder_jump : _GEN_54; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_56 = 4'h8 == io_ar_addr ? btb_8_pre_decoder_jump : _GEN_55; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_57 = 4'h9 == io_ar_addr ? btb_9_pre_decoder_jump : _GEN_56; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_58 = 4'ha == io_ar_addr ? btb_10_pre_decoder_jump : _GEN_57; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_59 = 4'hb == io_ar_addr ? btb_11_pre_decoder_jump : _GEN_58; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_60 = 4'hc == io_ar_addr ? btb_12_pre_decoder_jump : _GEN_59; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_61 = 4'hd == io_ar_addr ? btb_13_pre_decoder_jump : _GEN_60; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_62 = 4'he == io_ar_addr ? btb_14_pre_decoder_jump : _GEN_61; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_65 = 4'h1 == io_ar_addr ? btb_1_pre_decoder_branchD_flag : btb_0_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_66 = 4'h2 == io_ar_addr ? btb_2_pre_decoder_branchD_flag : _GEN_65; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_67 = 4'h3 == io_ar_addr ? btb_3_pre_decoder_branchD_flag : _GEN_66; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_68 = 4'h4 == io_ar_addr ? btb_4_pre_decoder_branchD_flag : _GEN_67; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_69 = 4'h5 == io_ar_addr ? btb_5_pre_decoder_branchD_flag : _GEN_68; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_70 = 4'h6 == io_ar_addr ? btb_6_pre_decoder_branchD_flag : _GEN_69; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_71 = 4'h7 == io_ar_addr ? btb_7_pre_decoder_branchD_flag : _GEN_70; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_72 = 4'h8 == io_ar_addr ? btb_8_pre_decoder_branchD_flag : _GEN_71; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_73 = 4'h9 == io_ar_addr ? btb_9_pre_decoder_branchD_flag : _GEN_72; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_74 = 4'ha == io_ar_addr ? btb_10_pre_decoder_branchD_flag : _GEN_73; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_75 = 4'hb == io_ar_addr ? btb_11_pre_decoder_branchD_flag : _GEN_74; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_76 = 4'hc == io_ar_addr ? btb_12_pre_decoder_branchD_flag : _GEN_75; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_77 = 4'hd == io_ar_addr ? btb_13_pre_decoder_branchD_flag : _GEN_76; // @[ports_lookup_table.scala 106:{12,12}]
  wire  _GEN_78 = 4'he == io_ar_addr ? btb_14_pre_decoder_branchD_flag : _GEN_77; // @[ports_lookup_table.scala 106:{12,12}]
  wire [7:0] _GEN_81 = 4'h1 == io_ar_addr ? btb_1_pre_lookup_value : btb_0_pre_lookup_value; // @[ports_lookup_table.scala 106:{12,12}]
  wire [7:0] _GEN_82 = 4'h2 == io_ar_addr ? btb_2_pre_lookup_value : _GEN_81; // @[ports_lookup_table.scala 106:{12,12}]
  wire [7:0] _GEN_83 = 4'h3 == io_ar_addr ? btb_3_pre_lookup_value : _GEN_82; // @[ports_lookup_table.scala 106:{12,12}]
  wire [7:0] _GEN_84 = 4'h4 == io_ar_addr ? btb_4_pre_lookup_value : _GEN_83; // @[ports_lookup_table.scala 106:{12,12}]
  wire [7:0] _GEN_85 = 4'h5 == io_ar_addr ? btb_5_pre_lookup_value : _GEN_84; // @[ports_lookup_table.scala 106:{12,12}]
  wire [7:0] _GEN_86 = 4'h6 == io_ar_addr ? btb_6_pre_lookup_value : _GEN_85; // @[ports_lookup_table.scala 106:{12,12}]
  wire [7:0] _GEN_87 = 4'h7 == io_ar_addr ? btb_7_pre_lookup_value : _GEN_86; // @[ports_lookup_table.scala 106:{12,12}]
  wire [7:0] _GEN_88 = 4'h8 == io_ar_addr ? btb_8_pre_lookup_value : _GEN_87; // @[ports_lookup_table.scala 106:{12,12}]
  wire [7:0] _GEN_89 = 4'h9 == io_ar_addr ? btb_9_pre_lookup_value : _GEN_88; // @[ports_lookup_table.scala 106:{12,12}]
  wire [7:0] _GEN_90 = 4'ha == io_ar_addr ? btb_10_pre_lookup_value : _GEN_89; // @[ports_lookup_table.scala 106:{12,12}]
  wire [7:0] _GEN_91 = 4'hb == io_ar_addr ? btb_11_pre_lookup_value : _GEN_90; // @[ports_lookup_table.scala 106:{12,12}]
  wire [7:0] _GEN_92 = 4'hc == io_ar_addr ? btb_12_pre_lookup_value : _GEN_91; // @[ports_lookup_table.scala 106:{12,12}]
  wire [7:0] _GEN_93 = 4'hd == io_ar_addr ? btb_13_pre_lookup_value : _GEN_92; // @[ports_lookup_table.scala 106:{12,12}]
  wire [7:0] _GEN_94 = 4'he == io_ar_addr ? btb_14_pre_lookup_value : _GEN_93; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_97 = 4'h1 == io_ar_addr ? btb_1_pre_bht : btb_0_pre_bht; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_98 = 4'h2 == io_ar_addr ? btb_2_pre_bht : _GEN_97; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_99 = 4'h3 == io_ar_addr ? btb_3_pre_bht : _GEN_98; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_100 = 4'h4 == io_ar_addr ? btb_4_pre_bht : _GEN_99; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_101 = 4'h5 == io_ar_addr ? btb_5_pre_bht : _GEN_100; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_102 = 4'h6 == io_ar_addr ? btb_6_pre_bht : _GEN_101; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_103 = 4'h7 == io_ar_addr ? btb_7_pre_bht : _GEN_102; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_104 = 4'h8 == io_ar_addr ? btb_8_pre_bht : _GEN_103; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_105 = 4'h9 == io_ar_addr ? btb_9_pre_bht : _GEN_104; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_106 = 4'ha == io_ar_addr ? btb_10_pre_bht : _GEN_105; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_107 = 4'hb == io_ar_addr ? btb_11_pre_bht : _GEN_106; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_108 = 4'hc == io_ar_addr ? btb_12_pre_bht : _GEN_107; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_109 = 4'hd == io_ar_addr ? btb_13_pre_bht : _GEN_108; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_110 = 4'he == io_ar_addr ? btb_14_pre_bht : _GEN_109; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_113 = 4'h1 == io_ar_addr ? btb_1_pre_pht : btb_0_pre_pht; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_114 = 4'h2 == io_ar_addr ? btb_2_pre_pht : _GEN_113; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_115 = 4'h3 == io_ar_addr ? btb_3_pre_pht : _GEN_114; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_116 = 4'h4 == io_ar_addr ? btb_4_pre_pht : _GEN_115; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_117 = 4'h5 == io_ar_addr ? btb_5_pre_pht : _GEN_116; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_118 = 4'h6 == io_ar_addr ? btb_6_pre_pht : _GEN_117; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_119 = 4'h7 == io_ar_addr ? btb_7_pre_pht : _GEN_118; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_120 = 4'h8 == io_ar_addr ? btb_8_pre_pht : _GEN_119; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_121 = 4'h9 == io_ar_addr ? btb_9_pre_pht : _GEN_120; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_122 = 4'ha == io_ar_addr ? btb_10_pre_pht : _GEN_121; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_123 = 4'hb == io_ar_addr ? btb_11_pre_pht : _GEN_122; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_124 = 4'hc == io_ar_addr ? btb_12_pre_pht : _GEN_123; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_125 = 4'hd == io_ar_addr ? btb_13_pre_pht : _GEN_124; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_126 = 4'he == io_ar_addr ? btb_14_pre_pht : _GEN_125; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_129 = 4'h1 == io_ar_addr ? btb_1_pre_hashcode : btb_0_pre_hashcode; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_130 = 4'h2 == io_ar_addr ? btb_2_pre_hashcode : _GEN_129; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_131 = 4'h3 == io_ar_addr ? btb_3_pre_hashcode : _GEN_130; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_132 = 4'h4 == io_ar_addr ? btb_4_pre_hashcode : _GEN_131; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_133 = 4'h5 == io_ar_addr ? btb_5_pre_hashcode : _GEN_132; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_134 = 4'h6 == io_ar_addr ? btb_6_pre_hashcode : _GEN_133; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_135 = 4'h7 == io_ar_addr ? btb_7_pre_hashcode : _GEN_134; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_136 = 4'h8 == io_ar_addr ? btb_8_pre_hashcode : _GEN_135; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_137 = 4'h9 == io_ar_addr ? btb_9_pre_hashcode : _GEN_136; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_138 = 4'ha == io_ar_addr ? btb_10_pre_hashcode : _GEN_137; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_139 = 4'hb == io_ar_addr ? btb_11_pre_hashcode : _GEN_138; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_140 = 4'hc == io_ar_addr ? btb_12_pre_hashcode : _GEN_139; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_141 = 4'hd == io_ar_addr ? btb_13_pre_hashcode : _GEN_140; // @[ports_lookup_table.scala 106:{12,12}]
  wire [3:0] _GEN_142 = 4'he == io_ar_addr ? btb_14_pre_hashcode : _GEN_141; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_145 = 4'h1 == io_ar_addr ? btb_1_pre_lookup_data : btb_0_pre_lookup_data; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_146 = 4'h2 == io_ar_addr ? btb_2_pre_lookup_data : _GEN_145; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_147 = 4'h3 == io_ar_addr ? btb_3_pre_lookup_data : _GEN_146; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_148 = 4'h4 == io_ar_addr ? btb_4_pre_lookup_data : _GEN_147; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_149 = 4'h5 == io_ar_addr ? btb_5_pre_lookup_data : _GEN_148; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_150 = 4'h6 == io_ar_addr ? btb_6_pre_lookup_data : _GEN_149; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_151 = 4'h7 == io_ar_addr ? btb_7_pre_lookup_data : _GEN_150; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_152 = 4'h8 == io_ar_addr ? btb_8_pre_lookup_data : _GEN_151; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_153 = 4'h9 == io_ar_addr ? btb_9_pre_lookup_data : _GEN_152; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_154 = 4'ha == io_ar_addr ? btb_10_pre_lookup_data : _GEN_153; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_155 = 4'hb == io_ar_addr ? btb_11_pre_lookup_data : _GEN_154; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_156 = 4'hc == io_ar_addr ? btb_12_pre_lookup_data : _GEN_155; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_157 = 4'hd == io_ar_addr ? btb_13_pre_lookup_data : _GEN_156; // @[ports_lookup_table.scala 106:{12,12}]
  wire [6:0] _GEN_158 = 4'he == io_ar_addr ? btb_14_pre_lookup_data : _GEN_157; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_161 = 4'h1 == io_ar_addr ? btb_1_pre_pc_target : btb_0_pre_pc_target; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_162 = 4'h2 == io_ar_addr ? btb_2_pre_pc_target : _GEN_161; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_163 = 4'h3 == io_ar_addr ? btb_3_pre_pc_target : _GEN_162; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_164 = 4'h4 == io_ar_addr ? btb_4_pre_pc_target : _GEN_163; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_165 = 4'h5 == io_ar_addr ? btb_5_pre_pc_target : _GEN_164; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_166 = 4'h6 == io_ar_addr ? btb_6_pre_pc_target : _GEN_165; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_167 = 4'h7 == io_ar_addr ? btb_7_pre_pc_target : _GEN_166; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_168 = 4'h8 == io_ar_addr ? btb_8_pre_pc_target : _GEN_167; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_169 = 4'h9 == io_ar_addr ? btb_9_pre_pc_target : _GEN_168; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_170 = 4'ha == io_ar_addr ? btb_10_pre_pc_target : _GEN_169; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_171 = 4'hb == io_ar_addr ? btb_11_pre_pc_target : _GEN_170; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_172 = 4'hc == io_ar_addr ? btb_12_pre_pc_target : _GEN_171; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_173 = 4'hd == io_ar_addr ? btb_13_pre_pc_target : _GEN_172; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_174 = 4'he == io_ar_addr ? btb_14_pre_pc_target : _GEN_173; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_177 = 4'h1 == io_ar_addr ? btb_1_exception_type : btb_0_exception_type; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_178 = 4'h2 == io_ar_addr ? btb_2_exception_type : _GEN_177; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_179 = 4'h3 == io_ar_addr ? btb_3_exception_type : _GEN_178; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_180 = 4'h4 == io_ar_addr ? btb_4_exception_type : _GEN_179; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_181 = 4'h5 == io_ar_addr ? btb_5_exception_type : _GEN_180; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_182 = 4'h6 == io_ar_addr ? btb_6_exception_type : _GEN_181; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_183 = 4'h7 == io_ar_addr ? btb_7_exception_type : _GEN_182; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_184 = 4'h8 == io_ar_addr ? btb_8_exception_type : _GEN_183; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_185 = 4'h9 == io_ar_addr ? btb_9_exception_type : _GEN_184; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_186 = 4'ha == io_ar_addr ? btb_10_exception_type : _GEN_185; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_187 = 4'hb == io_ar_addr ? btb_11_exception_type : _GEN_186; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_188 = 4'hc == io_ar_addr ? btb_12_exception_type : _GEN_187; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_189 = 4'hd == io_ar_addr ? btb_13_exception_type : _GEN_188; // @[ports_lookup_table.scala 106:{12,12}]
  wire [1:0] _GEN_190 = 4'he == io_ar_addr ? btb_14_exception_type : _GEN_189; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_193 = 4'h1 == io_ar_addr ? btb_1_inst : btb_0_inst; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_194 = 4'h2 == io_ar_addr ? btb_2_inst : _GEN_193; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_195 = 4'h3 == io_ar_addr ? btb_3_inst : _GEN_194; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_196 = 4'h4 == io_ar_addr ? btb_4_inst : _GEN_195; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_197 = 4'h5 == io_ar_addr ? btb_5_inst : _GEN_196; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_198 = 4'h6 == io_ar_addr ? btb_6_inst : _GEN_197; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_199 = 4'h7 == io_ar_addr ? btb_7_inst : _GEN_198; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_200 = 4'h8 == io_ar_addr ? btb_8_inst : _GEN_199; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_201 = 4'h9 == io_ar_addr ? btb_9_inst : _GEN_200; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_202 = 4'ha == io_ar_addr ? btb_10_inst : _GEN_201; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_203 = 4'hb == io_ar_addr ? btb_11_inst : _GEN_202; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_204 = 4'hc == io_ar_addr ? btb_12_inst : _GEN_203; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_205 = 4'hd == io_ar_addr ? btb_13_inst : _GEN_204; // @[ports_lookup_table.scala 106:{12,12}]
  wire [31:0] _GEN_206 = 4'he == io_ar_addr ? btb_14_inst : _GEN_205; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_209 = 4'h1 == io_ar_addr ? btb_1_pc : btb_0_pc; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_210 = 4'h2 == io_ar_addr ? btb_2_pc : _GEN_209; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_211 = 4'h3 == io_ar_addr ? btb_3_pc : _GEN_210; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_212 = 4'h4 == io_ar_addr ? btb_4_pc : _GEN_211; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_213 = 4'h5 == io_ar_addr ? btb_5_pc : _GEN_212; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_214 = 4'h6 == io_ar_addr ? btb_6_pc : _GEN_213; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_215 = 4'h7 == io_ar_addr ? btb_7_pc : _GEN_214; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_216 = 4'h8 == io_ar_addr ? btb_8_pc : _GEN_215; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_217 = 4'h9 == io_ar_addr ? btb_9_pc : _GEN_216; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_218 = 4'ha == io_ar_addr ? btb_10_pc : _GEN_217; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_219 = 4'hb == io_ar_addr ? btb_11_pc : _GEN_218; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_220 = 4'hc == io_ar_addr ? btb_12_pc : _GEN_219; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_221 = 4'hd == io_ar_addr ? btb_13_pc : _GEN_220; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_222 = 4'he == io_ar_addr ? btb_14_pc : _GEN_221; // @[ports_lookup_table.scala 106:{12,12}]
  wire [63:0] _GEN_238 = 4'h1 == io_aw_addr ? btb_1_pc : btb_0_pc; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_239 = 4'h1 == io_aw_addr ? btb_1_inst : btb_0_inst; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_240 = 4'h1 == io_aw_addr ? btb_1_exception_type : btb_0_exception_type; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_241 = 4'h1 == io_aw_addr ? btb_1_pre_pc_target : btb_0_pre_pc_target; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_242 = 4'h1 == io_aw_addr ? btb_1_pre_lookup_data : btb_0_pre_lookup_data; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_243 = 4'h1 == io_aw_addr ? btb_1_pre_hashcode : btb_0_pre_hashcode; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_244 = 4'h1 == io_aw_addr ? btb_1_pre_pht : btb_0_pre_pht; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_245 = 4'h1 == io_aw_addr ? btb_1_pre_bht : btb_0_pre_bht; // @[ports_lookup_table.scala 107:{27,27}]
  wire [7:0] _GEN_246 = 4'h1 == io_aw_addr ? btb_1_pre_lookup_value : btb_0_pre_lookup_value; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_247 = 4'h1 == io_aw_addr ? btb_1_pre_decoder_branchD_flag : btb_0_pre_decoder_branchD_flag; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_248 = 4'h1 == io_aw_addr ? btb_1_pre_decoder_jump : btb_0_pre_decoder_jump; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_249 = 4'h1 == io_aw_addr ? btb_1_pre_decoder_branchdata : btb_0_pre_decoder_branchdata; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_250 = 4'h1 == io_aw_addr ? btb_1_pre_decoder_jr : btb_0_pre_decoder_jr; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_251 = 4'h1 == io_aw_addr ? btb_1_true_branch_state : btb_0_true_branch_state; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_252 = 4'h2 == io_aw_addr ? btb_2_pc : _GEN_238; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_253 = 4'h2 == io_aw_addr ? btb_2_inst : _GEN_239; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_254 = 4'h2 == io_aw_addr ? btb_2_exception_type : _GEN_240; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_255 = 4'h2 == io_aw_addr ? btb_2_pre_pc_target : _GEN_241; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_256 = 4'h2 == io_aw_addr ? btb_2_pre_lookup_data : _GEN_242; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_257 = 4'h2 == io_aw_addr ? btb_2_pre_hashcode : _GEN_243; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_258 = 4'h2 == io_aw_addr ? btb_2_pre_pht : _GEN_244; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_259 = 4'h2 == io_aw_addr ? btb_2_pre_bht : _GEN_245; // @[ports_lookup_table.scala 107:{27,27}]
  wire [7:0] _GEN_260 = 4'h2 == io_aw_addr ? btb_2_pre_lookup_value : _GEN_246; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_261 = 4'h2 == io_aw_addr ? btb_2_pre_decoder_branchD_flag : _GEN_247; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_262 = 4'h2 == io_aw_addr ? btb_2_pre_decoder_jump : _GEN_248; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_263 = 4'h2 == io_aw_addr ? btb_2_pre_decoder_branchdata : _GEN_249; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_264 = 4'h2 == io_aw_addr ? btb_2_pre_decoder_jr : _GEN_250; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_265 = 4'h2 == io_aw_addr ? btb_2_true_branch_state : _GEN_251; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_266 = 4'h3 == io_aw_addr ? btb_3_pc : _GEN_252; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_267 = 4'h3 == io_aw_addr ? btb_3_inst : _GEN_253; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_268 = 4'h3 == io_aw_addr ? btb_3_exception_type : _GEN_254; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_269 = 4'h3 == io_aw_addr ? btb_3_pre_pc_target : _GEN_255; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_270 = 4'h3 == io_aw_addr ? btb_3_pre_lookup_data : _GEN_256; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_271 = 4'h3 == io_aw_addr ? btb_3_pre_hashcode : _GEN_257; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_272 = 4'h3 == io_aw_addr ? btb_3_pre_pht : _GEN_258; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_273 = 4'h3 == io_aw_addr ? btb_3_pre_bht : _GEN_259; // @[ports_lookup_table.scala 107:{27,27}]
  wire [7:0] _GEN_274 = 4'h3 == io_aw_addr ? btb_3_pre_lookup_value : _GEN_260; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_275 = 4'h3 == io_aw_addr ? btb_3_pre_decoder_branchD_flag : _GEN_261; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_276 = 4'h3 == io_aw_addr ? btb_3_pre_decoder_jump : _GEN_262; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_277 = 4'h3 == io_aw_addr ? btb_3_pre_decoder_branchdata : _GEN_263; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_278 = 4'h3 == io_aw_addr ? btb_3_pre_decoder_jr : _GEN_264; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_279 = 4'h3 == io_aw_addr ? btb_3_true_branch_state : _GEN_265; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_280 = 4'h4 == io_aw_addr ? btb_4_pc : _GEN_266; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_281 = 4'h4 == io_aw_addr ? btb_4_inst : _GEN_267; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_282 = 4'h4 == io_aw_addr ? btb_4_exception_type : _GEN_268; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_283 = 4'h4 == io_aw_addr ? btb_4_pre_pc_target : _GEN_269; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_284 = 4'h4 == io_aw_addr ? btb_4_pre_lookup_data : _GEN_270; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_285 = 4'h4 == io_aw_addr ? btb_4_pre_hashcode : _GEN_271; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_286 = 4'h4 == io_aw_addr ? btb_4_pre_pht : _GEN_272; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_287 = 4'h4 == io_aw_addr ? btb_4_pre_bht : _GEN_273; // @[ports_lookup_table.scala 107:{27,27}]
  wire [7:0] _GEN_288 = 4'h4 == io_aw_addr ? btb_4_pre_lookup_value : _GEN_274; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_289 = 4'h4 == io_aw_addr ? btb_4_pre_decoder_branchD_flag : _GEN_275; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_290 = 4'h4 == io_aw_addr ? btb_4_pre_decoder_jump : _GEN_276; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_291 = 4'h4 == io_aw_addr ? btb_4_pre_decoder_branchdata : _GEN_277; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_292 = 4'h4 == io_aw_addr ? btb_4_pre_decoder_jr : _GEN_278; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_293 = 4'h4 == io_aw_addr ? btb_4_true_branch_state : _GEN_279; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_294 = 4'h5 == io_aw_addr ? btb_5_pc : _GEN_280; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_295 = 4'h5 == io_aw_addr ? btb_5_inst : _GEN_281; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_296 = 4'h5 == io_aw_addr ? btb_5_exception_type : _GEN_282; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_297 = 4'h5 == io_aw_addr ? btb_5_pre_pc_target : _GEN_283; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_298 = 4'h5 == io_aw_addr ? btb_5_pre_lookup_data : _GEN_284; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_299 = 4'h5 == io_aw_addr ? btb_5_pre_hashcode : _GEN_285; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_300 = 4'h5 == io_aw_addr ? btb_5_pre_pht : _GEN_286; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_301 = 4'h5 == io_aw_addr ? btb_5_pre_bht : _GEN_287; // @[ports_lookup_table.scala 107:{27,27}]
  wire [7:0] _GEN_302 = 4'h5 == io_aw_addr ? btb_5_pre_lookup_value : _GEN_288; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_303 = 4'h5 == io_aw_addr ? btb_5_pre_decoder_branchD_flag : _GEN_289; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_304 = 4'h5 == io_aw_addr ? btb_5_pre_decoder_jump : _GEN_290; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_305 = 4'h5 == io_aw_addr ? btb_5_pre_decoder_branchdata : _GEN_291; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_306 = 4'h5 == io_aw_addr ? btb_5_pre_decoder_jr : _GEN_292; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_307 = 4'h5 == io_aw_addr ? btb_5_true_branch_state : _GEN_293; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_308 = 4'h6 == io_aw_addr ? btb_6_pc : _GEN_294; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_309 = 4'h6 == io_aw_addr ? btb_6_inst : _GEN_295; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_310 = 4'h6 == io_aw_addr ? btb_6_exception_type : _GEN_296; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_311 = 4'h6 == io_aw_addr ? btb_6_pre_pc_target : _GEN_297; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_312 = 4'h6 == io_aw_addr ? btb_6_pre_lookup_data : _GEN_298; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_313 = 4'h6 == io_aw_addr ? btb_6_pre_hashcode : _GEN_299; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_314 = 4'h6 == io_aw_addr ? btb_6_pre_pht : _GEN_300; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_315 = 4'h6 == io_aw_addr ? btb_6_pre_bht : _GEN_301; // @[ports_lookup_table.scala 107:{27,27}]
  wire [7:0] _GEN_316 = 4'h6 == io_aw_addr ? btb_6_pre_lookup_value : _GEN_302; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_317 = 4'h6 == io_aw_addr ? btb_6_pre_decoder_branchD_flag : _GEN_303; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_318 = 4'h6 == io_aw_addr ? btb_6_pre_decoder_jump : _GEN_304; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_319 = 4'h6 == io_aw_addr ? btb_6_pre_decoder_branchdata : _GEN_305; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_320 = 4'h6 == io_aw_addr ? btb_6_pre_decoder_jr : _GEN_306; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_321 = 4'h6 == io_aw_addr ? btb_6_true_branch_state : _GEN_307; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_322 = 4'h7 == io_aw_addr ? btb_7_pc : _GEN_308; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_323 = 4'h7 == io_aw_addr ? btb_7_inst : _GEN_309; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_324 = 4'h7 == io_aw_addr ? btb_7_exception_type : _GEN_310; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_325 = 4'h7 == io_aw_addr ? btb_7_pre_pc_target : _GEN_311; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_326 = 4'h7 == io_aw_addr ? btb_7_pre_lookup_data : _GEN_312; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_327 = 4'h7 == io_aw_addr ? btb_7_pre_hashcode : _GEN_313; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_328 = 4'h7 == io_aw_addr ? btb_7_pre_pht : _GEN_314; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_329 = 4'h7 == io_aw_addr ? btb_7_pre_bht : _GEN_315; // @[ports_lookup_table.scala 107:{27,27}]
  wire [7:0] _GEN_330 = 4'h7 == io_aw_addr ? btb_7_pre_lookup_value : _GEN_316; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_331 = 4'h7 == io_aw_addr ? btb_7_pre_decoder_branchD_flag : _GEN_317; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_332 = 4'h7 == io_aw_addr ? btb_7_pre_decoder_jump : _GEN_318; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_333 = 4'h7 == io_aw_addr ? btb_7_pre_decoder_branchdata : _GEN_319; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_334 = 4'h7 == io_aw_addr ? btb_7_pre_decoder_jr : _GEN_320; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_335 = 4'h7 == io_aw_addr ? btb_7_true_branch_state : _GEN_321; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_336 = 4'h8 == io_aw_addr ? btb_8_pc : _GEN_322; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_337 = 4'h8 == io_aw_addr ? btb_8_inst : _GEN_323; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_338 = 4'h8 == io_aw_addr ? btb_8_exception_type : _GEN_324; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_339 = 4'h8 == io_aw_addr ? btb_8_pre_pc_target : _GEN_325; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_340 = 4'h8 == io_aw_addr ? btb_8_pre_lookup_data : _GEN_326; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_341 = 4'h8 == io_aw_addr ? btb_8_pre_hashcode : _GEN_327; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_342 = 4'h8 == io_aw_addr ? btb_8_pre_pht : _GEN_328; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_343 = 4'h8 == io_aw_addr ? btb_8_pre_bht : _GEN_329; // @[ports_lookup_table.scala 107:{27,27}]
  wire [7:0] _GEN_344 = 4'h8 == io_aw_addr ? btb_8_pre_lookup_value : _GEN_330; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_345 = 4'h8 == io_aw_addr ? btb_8_pre_decoder_branchD_flag : _GEN_331; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_346 = 4'h8 == io_aw_addr ? btb_8_pre_decoder_jump : _GEN_332; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_347 = 4'h8 == io_aw_addr ? btb_8_pre_decoder_branchdata : _GEN_333; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_348 = 4'h8 == io_aw_addr ? btb_8_pre_decoder_jr : _GEN_334; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_349 = 4'h8 == io_aw_addr ? btb_8_true_branch_state : _GEN_335; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_350 = 4'h9 == io_aw_addr ? btb_9_pc : _GEN_336; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_351 = 4'h9 == io_aw_addr ? btb_9_inst : _GEN_337; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_352 = 4'h9 == io_aw_addr ? btb_9_exception_type : _GEN_338; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_353 = 4'h9 == io_aw_addr ? btb_9_pre_pc_target : _GEN_339; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_354 = 4'h9 == io_aw_addr ? btb_9_pre_lookup_data : _GEN_340; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_355 = 4'h9 == io_aw_addr ? btb_9_pre_hashcode : _GEN_341; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_356 = 4'h9 == io_aw_addr ? btb_9_pre_pht : _GEN_342; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_357 = 4'h9 == io_aw_addr ? btb_9_pre_bht : _GEN_343; // @[ports_lookup_table.scala 107:{27,27}]
  wire [7:0] _GEN_358 = 4'h9 == io_aw_addr ? btb_9_pre_lookup_value : _GEN_344; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_359 = 4'h9 == io_aw_addr ? btb_9_pre_decoder_branchD_flag : _GEN_345; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_360 = 4'h9 == io_aw_addr ? btb_9_pre_decoder_jump : _GEN_346; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_361 = 4'h9 == io_aw_addr ? btb_9_pre_decoder_branchdata : _GEN_347; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_362 = 4'h9 == io_aw_addr ? btb_9_pre_decoder_jr : _GEN_348; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_363 = 4'h9 == io_aw_addr ? btb_9_true_branch_state : _GEN_349; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_364 = 4'ha == io_aw_addr ? btb_10_pc : _GEN_350; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_365 = 4'ha == io_aw_addr ? btb_10_inst : _GEN_351; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_366 = 4'ha == io_aw_addr ? btb_10_exception_type : _GEN_352; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_367 = 4'ha == io_aw_addr ? btb_10_pre_pc_target : _GEN_353; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_368 = 4'ha == io_aw_addr ? btb_10_pre_lookup_data : _GEN_354; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_369 = 4'ha == io_aw_addr ? btb_10_pre_hashcode : _GEN_355; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_370 = 4'ha == io_aw_addr ? btb_10_pre_pht : _GEN_356; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_371 = 4'ha == io_aw_addr ? btb_10_pre_bht : _GEN_357; // @[ports_lookup_table.scala 107:{27,27}]
  wire [7:0] _GEN_372 = 4'ha == io_aw_addr ? btb_10_pre_lookup_value : _GEN_358; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_373 = 4'ha == io_aw_addr ? btb_10_pre_decoder_branchD_flag : _GEN_359; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_374 = 4'ha == io_aw_addr ? btb_10_pre_decoder_jump : _GEN_360; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_375 = 4'ha == io_aw_addr ? btb_10_pre_decoder_branchdata : _GEN_361; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_376 = 4'ha == io_aw_addr ? btb_10_pre_decoder_jr : _GEN_362; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_377 = 4'ha == io_aw_addr ? btb_10_true_branch_state : _GEN_363; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_378 = 4'hb == io_aw_addr ? btb_11_pc : _GEN_364; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_379 = 4'hb == io_aw_addr ? btb_11_inst : _GEN_365; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_380 = 4'hb == io_aw_addr ? btb_11_exception_type : _GEN_366; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_381 = 4'hb == io_aw_addr ? btb_11_pre_pc_target : _GEN_367; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_382 = 4'hb == io_aw_addr ? btb_11_pre_lookup_data : _GEN_368; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_383 = 4'hb == io_aw_addr ? btb_11_pre_hashcode : _GEN_369; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_384 = 4'hb == io_aw_addr ? btb_11_pre_pht : _GEN_370; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_385 = 4'hb == io_aw_addr ? btb_11_pre_bht : _GEN_371; // @[ports_lookup_table.scala 107:{27,27}]
  wire [7:0] _GEN_386 = 4'hb == io_aw_addr ? btb_11_pre_lookup_value : _GEN_372; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_387 = 4'hb == io_aw_addr ? btb_11_pre_decoder_branchD_flag : _GEN_373; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_388 = 4'hb == io_aw_addr ? btb_11_pre_decoder_jump : _GEN_374; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_389 = 4'hb == io_aw_addr ? btb_11_pre_decoder_branchdata : _GEN_375; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_390 = 4'hb == io_aw_addr ? btb_11_pre_decoder_jr : _GEN_376; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_391 = 4'hb == io_aw_addr ? btb_11_true_branch_state : _GEN_377; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_392 = 4'hc == io_aw_addr ? btb_12_pc : _GEN_378; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_393 = 4'hc == io_aw_addr ? btb_12_inst : _GEN_379; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_394 = 4'hc == io_aw_addr ? btb_12_exception_type : _GEN_380; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_395 = 4'hc == io_aw_addr ? btb_12_pre_pc_target : _GEN_381; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_396 = 4'hc == io_aw_addr ? btb_12_pre_lookup_data : _GEN_382; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_397 = 4'hc == io_aw_addr ? btb_12_pre_hashcode : _GEN_383; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_398 = 4'hc == io_aw_addr ? btb_12_pre_pht : _GEN_384; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_399 = 4'hc == io_aw_addr ? btb_12_pre_bht : _GEN_385; // @[ports_lookup_table.scala 107:{27,27}]
  wire [7:0] _GEN_400 = 4'hc == io_aw_addr ? btb_12_pre_lookup_value : _GEN_386; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_401 = 4'hc == io_aw_addr ? btb_12_pre_decoder_branchD_flag : _GEN_387; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_402 = 4'hc == io_aw_addr ? btb_12_pre_decoder_jump : _GEN_388; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_403 = 4'hc == io_aw_addr ? btb_12_pre_decoder_branchdata : _GEN_389; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_404 = 4'hc == io_aw_addr ? btb_12_pre_decoder_jr : _GEN_390; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_405 = 4'hc == io_aw_addr ? btb_12_true_branch_state : _GEN_391; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_406 = 4'hd == io_aw_addr ? btb_13_pc : _GEN_392; // @[ports_lookup_table.scala 107:{27,27}]
  wire [31:0] _GEN_407 = 4'hd == io_aw_addr ? btb_13_inst : _GEN_393; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_408 = 4'hd == io_aw_addr ? btb_13_exception_type : _GEN_394; // @[ports_lookup_table.scala 107:{27,27}]
  wire [63:0] _GEN_409 = 4'hd == io_aw_addr ? btb_13_pre_pc_target : _GEN_395; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_410 = 4'hd == io_aw_addr ? btb_13_pre_lookup_data : _GEN_396; // @[ports_lookup_table.scala 107:{27,27}]
  wire [3:0] _GEN_411 = 4'hd == io_aw_addr ? btb_13_pre_hashcode : _GEN_397; // @[ports_lookup_table.scala 107:{27,27}]
  wire [1:0] _GEN_412 = 4'hd == io_aw_addr ? btb_13_pre_pht : _GEN_398; // @[ports_lookup_table.scala 107:{27,27}]
  wire [6:0] _GEN_413 = 4'hd == io_aw_addr ? btb_13_pre_bht : _GEN_399; // @[ports_lookup_table.scala 107:{27,27}]
  wire [7:0] _GEN_414 = 4'hd == io_aw_addr ? btb_13_pre_lookup_value : _GEN_400; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_415 = 4'hd == io_aw_addr ? btb_13_pre_decoder_branchD_flag : _GEN_401; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_416 = 4'hd == io_aw_addr ? btb_13_pre_decoder_jump : _GEN_402; // @[ports_lookup_table.scala 107:{27,27}]
  wire [5:0] _GEN_417 = 4'hd == io_aw_addr ? btb_13_pre_decoder_branchdata : _GEN_403; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_418 = 4'hd == io_aw_addr ? btb_13_pre_decoder_jr : _GEN_404; // @[ports_lookup_table.scala 107:{27,27}]
  wire  _GEN_419 = 4'hd == io_aw_addr ? btb_13_true_branch_state : _GEN_405; // @[ports_lookup_table.scala 107:{27,27}]
  assign io_out_pc = 4'hf == io_ar_addr ? btb_15_pc : _GEN_222; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_inst = 4'hf == io_ar_addr ? btb_15_inst : _GEN_206; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_exception_type = 4'hf == io_ar_addr ? btb_15_exception_type : _GEN_190; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_pre_pc_target = 4'hf == io_ar_addr ? btb_15_pre_pc_target : _GEN_174; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_pre_lookup_data = 4'hf == io_ar_addr ? btb_15_pre_lookup_data : _GEN_158; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_pre_hashcode = 4'hf == io_ar_addr ? btb_15_pre_hashcode : _GEN_142; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_pre_pht = 4'hf == io_ar_addr ? btb_15_pre_pht : _GEN_126; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_pre_bht = 4'hf == io_ar_addr ? btb_15_pre_bht : _GEN_110; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_pre_lookup_value = 4'hf == io_ar_addr ? btb_15_pre_lookup_value : _GEN_94; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_pre_decoder_branchD_flag = 4'hf == io_ar_addr ? btb_15_pre_decoder_branchD_flag : _GEN_78; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_pre_decoder_jump = 4'hf == io_ar_addr ? btb_15_pre_decoder_jump : _GEN_62; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_pre_decoder_branchdata = 4'hf == io_ar_addr ? btb_15_pre_decoder_branchdata : _GEN_46; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_pre_decoder_jr = 4'hf == io_ar_addr ? btb_15_pre_decoder_jr : _GEN_30; // @[ports_lookup_table.scala 106:{12,12}]
  assign io_out_true_branch_state = 4'hf == io_ar_addr ? btb_15_true_branch_state : _GEN_14; // @[ports_lookup_table.scala 106:{12,12}]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_0_pc <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_0_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin
        btb_0_pc <= btb_15_pc;
      end else if (4'he == io_aw_addr) begin
        btb_0_pc <= btb_14_pc;
      end else begin
        btb_0_pc <= _GEN_406;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_0_inst <= 32'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_0_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin
        btb_0_inst <= btb_15_inst;
      end else if (4'he == io_aw_addr) begin
        btb_0_inst <= btb_14_inst;
      end else begin
        btb_0_inst <= _GEN_407;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_0_exception_type <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_0_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin
        btb_0_exception_type <= btb_15_exception_type;
      end else if (4'he == io_aw_addr) begin
        btb_0_exception_type <= btb_14_exception_type;
      end else begin
        btb_0_exception_type <= _GEN_408;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_0_pre_pc_target <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_0_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin
        btb_0_pre_pc_target <= btb_15_pre_pc_target;
      end else if (4'he == io_aw_addr) begin
        btb_0_pre_pc_target <= btb_14_pre_pc_target;
      end else begin
        btb_0_pre_pc_target <= _GEN_409;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_0_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_0_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin
        btb_0_pre_lookup_data <= btb_15_pre_lookup_data;
      end else if (4'he == io_aw_addr) begin
        btb_0_pre_lookup_data <= btb_14_pre_lookup_data;
      end else begin
        btb_0_pre_lookup_data <= _GEN_410;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_0_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_0_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin
        btb_0_pre_hashcode <= btb_15_pre_hashcode;
      end else if (4'he == io_aw_addr) begin
        btb_0_pre_hashcode <= btb_14_pre_hashcode;
      end else begin
        btb_0_pre_hashcode <= _GEN_411;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_0_pre_pht <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_0_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin
        btb_0_pre_pht <= btb_15_pre_pht;
      end else if (4'he == io_aw_addr) begin
        btb_0_pre_pht <= btb_14_pre_pht;
      end else begin
        btb_0_pre_pht <= _GEN_412;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_0_pre_bht <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_0_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin
        btb_0_pre_bht <= btb_15_pre_bht;
      end else if (4'he == io_aw_addr) begin
        btb_0_pre_bht <= btb_14_pre_bht;
      end else begin
        btb_0_pre_bht <= _GEN_413;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_0_pre_lookup_value <= 8'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_0_pre_lookup_value <= io_in_pre_lookup_value;
      end else if (4'hf == io_aw_addr) begin
        btb_0_pre_lookup_value <= btb_15_pre_lookup_value;
      end else if (4'he == io_aw_addr) begin
        btb_0_pre_lookup_value <= btb_14_pre_lookup_value;
      end else begin
        btb_0_pre_lookup_value <= _GEN_414;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_0_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_0_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin
        btb_0_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag;
      end else if (4'he == io_aw_addr) begin
        btb_0_pre_decoder_branchD_flag <= btb_14_pre_decoder_branchD_flag;
      end else begin
        btb_0_pre_decoder_branchD_flag <= _GEN_415;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_0_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_0_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin
        btb_0_pre_decoder_jump <= btb_15_pre_decoder_jump;
      end else if (4'he == io_aw_addr) begin
        btb_0_pre_decoder_jump <= btb_14_pre_decoder_jump;
      end else begin
        btb_0_pre_decoder_jump <= _GEN_416;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_0_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_0_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin
        btb_0_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata;
      end else if (4'he == io_aw_addr) begin
        btb_0_pre_decoder_branchdata <= btb_14_pre_decoder_branchdata;
      end else begin
        btb_0_pre_decoder_branchdata <= _GEN_417;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_0_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_0_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin
        btb_0_pre_decoder_jr <= btb_15_pre_decoder_jr;
      end else if (4'he == io_aw_addr) begin
        btb_0_pre_decoder_jr <= btb_14_pre_decoder_jr;
      end else begin
        btb_0_pre_decoder_jr <= _GEN_418;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_0_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_0_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin
        btb_0_true_branch_state <= btb_15_true_branch_state;
      end else if (4'he == io_aw_addr) begin
        btb_0_true_branch_state <= btb_14_true_branch_state;
      end else begin
        btb_0_true_branch_state <= _GEN_419;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_1_pc <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_1_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin
        btb_1_pc <= btb_15_pc;
      end else if (4'he == io_aw_addr) begin
        btb_1_pc <= btb_14_pc;
      end else begin
        btb_1_pc <= _GEN_406;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_1_inst <= 32'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_1_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin
        btb_1_inst <= btb_15_inst;
      end else if (4'he == io_aw_addr) begin
        btb_1_inst <= btb_14_inst;
      end else begin
        btb_1_inst <= _GEN_407;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_1_exception_type <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_1_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin
        btb_1_exception_type <= btb_15_exception_type;
      end else if (4'he == io_aw_addr) begin
        btb_1_exception_type <= btb_14_exception_type;
      end else begin
        btb_1_exception_type <= _GEN_408;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_1_pre_pc_target <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_1_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin
        btb_1_pre_pc_target <= btb_15_pre_pc_target;
      end else if (4'he == io_aw_addr) begin
        btb_1_pre_pc_target <= btb_14_pre_pc_target;
      end else begin
        btb_1_pre_pc_target <= _GEN_409;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_1_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_1_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin
        btb_1_pre_lookup_data <= btb_15_pre_lookup_data;
      end else if (4'he == io_aw_addr) begin
        btb_1_pre_lookup_data <= btb_14_pre_lookup_data;
      end else begin
        btb_1_pre_lookup_data <= _GEN_410;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_1_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_1_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin
        btb_1_pre_hashcode <= btb_15_pre_hashcode;
      end else if (4'he == io_aw_addr) begin
        btb_1_pre_hashcode <= btb_14_pre_hashcode;
      end else begin
        btb_1_pre_hashcode <= _GEN_411;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_1_pre_pht <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_1_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin
        btb_1_pre_pht <= btb_15_pre_pht;
      end else if (4'he == io_aw_addr) begin
        btb_1_pre_pht <= btb_14_pre_pht;
      end else begin
        btb_1_pre_pht <= _GEN_412;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_1_pre_bht <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_1_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin
        btb_1_pre_bht <= btb_15_pre_bht;
      end else if (4'he == io_aw_addr) begin
        btb_1_pre_bht <= btb_14_pre_bht;
      end else begin
        btb_1_pre_bht <= _GEN_413;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_1_pre_lookup_value <= 8'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_1_pre_lookup_value <= io_in_pre_lookup_value;
      end else if (4'hf == io_aw_addr) begin
        btb_1_pre_lookup_value <= btb_15_pre_lookup_value;
      end else if (4'he == io_aw_addr) begin
        btb_1_pre_lookup_value <= btb_14_pre_lookup_value;
      end else begin
        btb_1_pre_lookup_value <= _GEN_414;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_1_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_1_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin
        btb_1_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag;
      end else if (4'he == io_aw_addr) begin
        btb_1_pre_decoder_branchD_flag <= btb_14_pre_decoder_branchD_flag;
      end else begin
        btb_1_pre_decoder_branchD_flag <= _GEN_415;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_1_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_1_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin
        btb_1_pre_decoder_jump <= btb_15_pre_decoder_jump;
      end else if (4'he == io_aw_addr) begin
        btb_1_pre_decoder_jump <= btb_14_pre_decoder_jump;
      end else begin
        btb_1_pre_decoder_jump <= _GEN_416;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_1_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_1_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin
        btb_1_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata;
      end else if (4'he == io_aw_addr) begin
        btb_1_pre_decoder_branchdata <= btb_14_pre_decoder_branchdata;
      end else begin
        btb_1_pre_decoder_branchdata <= _GEN_417;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_1_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_1_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin
        btb_1_pre_decoder_jr <= btb_15_pre_decoder_jr;
      end else if (4'he == io_aw_addr) begin
        btb_1_pre_decoder_jr <= btb_14_pre_decoder_jr;
      end else begin
        btb_1_pre_decoder_jr <= _GEN_418;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_1_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_1_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin
        btb_1_true_branch_state <= btb_15_true_branch_state;
      end else if (4'he == io_aw_addr) begin
        btb_1_true_branch_state <= btb_14_true_branch_state;
      end else begin
        btb_1_true_branch_state <= _GEN_419;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_2_pc <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_2_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin
        btb_2_pc <= btb_15_pc;
      end else if (4'he == io_aw_addr) begin
        btb_2_pc <= btb_14_pc;
      end else begin
        btb_2_pc <= _GEN_406;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_2_inst <= 32'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_2_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin
        btb_2_inst <= btb_15_inst;
      end else if (4'he == io_aw_addr) begin
        btb_2_inst <= btb_14_inst;
      end else begin
        btb_2_inst <= _GEN_407;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_2_exception_type <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_2_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin
        btb_2_exception_type <= btb_15_exception_type;
      end else if (4'he == io_aw_addr) begin
        btb_2_exception_type <= btb_14_exception_type;
      end else begin
        btb_2_exception_type <= _GEN_408;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_2_pre_pc_target <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_2_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin
        btb_2_pre_pc_target <= btb_15_pre_pc_target;
      end else if (4'he == io_aw_addr) begin
        btb_2_pre_pc_target <= btb_14_pre_pc_target;
      end else begin
        btb_2_pre_pc_target <= _GEN_409;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_2_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_2_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin
        btb_2_pre_lookup_data <= btb_15_pre_lookup_data;
      end else if (4'he == io_aw_addr) begin
        btb_2_pre_lookup_data <= btb_14_pre_lookup_data;
      end else begin
        btb_2_pre_lookup_data <= _GEN_410;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_2_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_2_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin
        btb_2_pre_hashcode <= btb_15_pre_hashcode;
      end else if (4'he == io_aw_addr) begin
        btb_2_pre_hashcode <= btb_14_pre_hashcode;
      end else begin
        btb_2_pre_hashcode <= _GEN_411;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_2_pre_pht <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_2_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin
        btb_2_pre_pht <= btb_15_pre_pht;
      end else if (4'he == io_aw_addr) begin
        btb_2_pre_pht <= btb_14_pre_pht;
      end else begin
        btb_2_pre_pht <= _GEN_412;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_2_pre_bht <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_2_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin
        btb_2_pre_bht <= btb_15_pre_bht;
      end else if (4'he == io_aw_addr) begin
        btb_2_pre_bht <= btb_14_pre_bht;
      end else begin
        btb_2_pre_bht <= _GEN_413;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_2_pre_lookup_value <= 8'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_2_pre_lookup_value <= io_in_pre_lookup_value;
      end else if (4'hf == io_aw_addr) begin
        btb_2_pre_lookup_value <= btb_15_pre_lookup_value;
      end else if (4'he == io_aw_addr) begin
        btb_2_pre_lookup_value <= btb_14_pre_lookup_value;
      end else begin
        btb_2_pre_lookup_value <= _GEN_414;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_2_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_2_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin
        btb_2_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag;
      end else if (4'he == io_aw_addr) begin
        btb_2_pre_decoder_branchD_flag <= btb_14_pre_decoder_branchD_flag;
      end else begin
        btb_2_pre_decoder_branchD_flag <= _GEN_415;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_2_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_2_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin
        btb_2_pre_decoder_jump <= btb_15_pre_decoder_jump;
      end else if (4'he == io_aw_addr) begin
        btb_2_pre_decoder_jump <= btb_14_pre_decoder_jump;
      end else begin
        btb_2_pre_decoder_jump <= _GEN_416;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_2_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_2_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin
        btb_2_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata;
      end else if (4'he == io_aw_addr) begin
        btb_2_pre_decoder_branchdata <= btb_14_pre_decoder_branchdata;
      end else begin
        btb_2_pre_decoder_branchdata <= _GEN_417;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_2_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_2_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin
        btb_2_pre_decoder_jr <= btb_15_pre_decoder_jr;
      end else if (4'he == io_aw_addr) begin
        btb_2_pre_decoder_jr <= btb_14_pre_decoder_jr;
      end else begin
        btb_2_pre_decoder_jr <= _GEN_418;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_2_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_2_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin
        btb_2_true_branch_state <= btb_15_true_branch_state;
      end else if (4'he == io_aw_addr) begin
        btb_2_true_branch_state <= btb_14_true_branch_state;
      end else begin
        btb_2_true_branch_state <= _GEN_419;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_3_pc <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_3_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin
        btb_3_pc <= btb_15_pc;
      end else if (4'he == io_aw_addr) begin
        btb_3_pc <= btb_14_pc;
      end else begin
        btb_3_pc <= _GEN_406;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_3_inst <= 32'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_3_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin
        btb_3_inst <= btb_15_inst;
      end else if (4'he == io_aw_addr) begin
        btb_3_inst <= btb_14_inst;
      end else begin
        btb_3_inst <= _GEN_407;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_3_exception_type <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_3_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin
        btb_3_exception_type <= btb_15_exception_type;
      end else if (4'he == io_aw_addr) begin
        btb_3_exception_type <= btb_14_exception_type;
      end else begin
        btb_3_exception_type <= _GEN_408;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_3_pre_pc_target <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_3_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin
        btb_3_pre_pc_target <= btb_15_pre_pc_target;
      end else if (4'he == io_aw_addr) begin
        btb_3_pre_pc_target <= btb_14_pre_pc_target;
      end else begin
        btb_3_pre_pc_target <= _GEN_409;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_3_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_3_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin
        btb_3_pre_lookup_data <= btb_15_pre_lookup_data;
      end else if (4'he == io_aw_addr) begin
        btb_3_pre_lookup_data <= btb_14_pre_lookup_data;
      end else begin
        btb_3_pre_lookup_data <= _GEN_410;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_3_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_3_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin
        btb_3_pre_hashcode <= btb_15_pre_hashcode;
      end else if (4'he == io_aw_addr) begin
        btb_3_pre_hashcode <= btb_14_pre_hashcode;
      end else begin
        btb_3_pre_hashcode <= _GEN_411;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_3_pre_pht <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_3_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin
        btb_3_pre_pht <= btb_15_pre_pht;
      end else if (4'he == io_aw_addr) begin
        btb_3_pre_pht <= btb_14_pre_pht;
      end else begin
        btb_3_pre_pht <= _GEN_412;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_3_pre_bht <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_3_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin
        btb_3_pre_bht <= btb_15_pre_bht;
      end else if (4'he == io_aw_addr) begin
        btb_3_pre_bht <= btb_14_pre_bht;
      end else begin
        btb_3_pre_bht <= _GEN_413;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_3_pre_lookup_value <= 8'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_3_pre_lookup_value <= io_in_pre_lookup_value;
      end else if (4'hf == io_aw_addr) begin
        btb_3_pre_lookup_value <= btb_15_pre_lookup_value;
      end else if (4'he == io_aw_addr) begin
        btb_3_pre_lookup_value <= btb_14_pre_lookup_value;
      end else begin
        btb_3_pre_lookup_value <= _GEN_414;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_3_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_3_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin
        btb_3_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag;
      end else if (4'he == io_aw_addr) begin
        btb_3_pre_decoder_branchD_flag <= btb_14_pre_decoder_branchD_flag;
      end else begin
        btb_3_pre_decoder_branchD_flag <= _GEN_415;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_3_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_3_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin
        btb_3_pre_decoder_jump <= btb_15_pre_decoder_jump;
      end else if (4'he == io_aw_addr) begin
        btb_3_pre_decoder_jump <= btb_14_pre_decoder_jump;
      end else begin
        btb_3_pre_decoder_jump <= _GEN_416;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_3_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_3_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin
        btb_3_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata;
      end else if (4'he == io_aw_addr) begin
        btb_3_pre_decoder_branchdata <= btb_14_pre_decoder_branchdata;
      end else begin
        btb_3_pre_decoder_branchdata <= _GEN_417;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_3_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_3_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin
        btb_3_pre_decoder_jr <= btb_15_pre_decoder_jr;
      end else if (4'he == io_aw_addr) begin
        btb_3_pre_decoder_jr <= btb_14_pre_decoder_jr;
      end else begin
        btb_3_pre_decoder_jr <= _GEN_418;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_3_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_3_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin
        btb_3_true_branch_state <= btb_15_true_branch_state;
      end else if (4'he == io_aw_addr) begin
        btb_3_true_branch_state <= btb_14_true_branch_state;
      end else begin
        btb_3_true_branch_state <= _GEN_419;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_4_pc <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_4_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin
        btb_4_pc <= btb_15_pc;
      end else if (4'he == io_aw_addr) begin
        btb_4_pc <= btb_14_pc;
      end else begin
        btb_4_pc <= _GEN_406;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_4_inst <= 32'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_4_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin
        btb_4_inst <= btb_15_inst;
      end else if (4'he == io_aw_addr) begin
        btb_4_inst <= btb_14_inst;
      end else begin
        btb_4_inst <= _GEN_407;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_4_exception_type <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_4_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin
        btb_4_exception_type <= btb_15_exception_type;
      end else if (4'he == io_aw_addr) begin
        btb_4_exception_type <= btb_14_exception_type;
      end else begin
        btb_4_exception_type <= _GEN_408;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_4_pre_pc_target <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_4_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin
        btb_4_pre_pc_target <= btb_15_pre_pc_target;
      end else if (4'he == io_aw_addr) begin
        btb_4_pre_pc_target <= btb_14_pre_pc_target;
      end else begin
        btb_4_pre_pc_target <= _GEN_409;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_4_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_4_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin
        btb_4_pre_lookup_data <= btb_15_pre_lookup_data;
      end else if (4'he == io_aw_addr) begin
        btb_4_pre_lookup_data <= btb_14_pre_lookup_data;
      end else begin
        btb_4_pre_lookup_data <= _GEN_410;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_4_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_4_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin
        btb_4_pre_hashcode <= btb_15_pre_hashcode;
      end else if (4'he == io_aw_addr) begin
        btb_4_pre_hashcode <= btb_14_pre_hashcode;
      end else begin
        btb_4_pre_hashcode <= _GEN_411;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_4_pre_pht <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_4_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin
        btb_4_pre_pht <= btb_15_pre_pht;
      end else if (4'he == io_aw_addr) begin
        btb_4_pre_pht <= btb_14_pre_pht;
      end else begin
        btb_4_pre_pht <= _GEN_412;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_4_pre_bht <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_4_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin
        btb_4_pre_bht <= btb_15_pre_bht;
      end else if (4'he == io_aw_addr) begin
        btb_4_pre_bht <= btb_14_pre_bht;
      end else begin
        btb_4_pre_bht <= _GEN_413;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_4_pre_lookup_value <= 8'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_4_pre_lookup_value <= io_in_pre_lookup_value;
      end else if (4'hf == io_aw_addr) begin
        btb_4_pre_lookup_value <= btb_15_pre_lookup_value;
      end else if (4'he == io_aw_addr) begin
        btb_4_pre_lookup_value <= btb_14_pre_lookup_value;
      end else begin
        btb_4_pre_lookup_value <= _GEN_414;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_4_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_4_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin
        btb_4_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag;
      end else if (4'he == io_aw_addr) begin
        btb_4_pre_decoder_branchD_flag <= btb_14_pre_decoder_branchD_flag;
      end else begin
        btb_4_pre_decoder_branchD_flag <= _GEN_415;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_4_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_4_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin
        btb_4_pre_decoder_jump <= btb_15_pre_decoder_jump;
      end else if (4'he == io_aw_addr) begin
        btb_4_pre_decoder_jump <= btb_14_pre_decoder_jump;
      end else begin
        btb_4_pre_decoder_jump <= _GEN_416;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_4_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_4_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin
        btb_4_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata;
      end else if (4'he == io_aw_addr) begin
        btb_4_pre_decoder_branchdata <= btb_14_pre_decoder_branchdata;
      end else begin
        btb_4_pre_decoder_branchdata <= _GEN_417;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_4_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_4_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin
        btb_4_pre_decoder_jr <= btb_15_pre_decoder_jr;
      end else if (4'he == io_aw_addr) begin
        btb_4_pre_decoder_jr <= btb_14_pre_decoder_jr;
      end else begin
        btb_4_pre_decoder_jr <= _GEN_418;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_4_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_4_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin
        btb_4_true_branch_state <= btb_15_true_branch_state;
      end else if (4'he == io_aw_addr) begin
        btb_4_true_branch_state <= btb_14_true_branch_state;
      end else begin
        btb_4_true_branch_state <= _GEN_419;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_5_pc <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_5_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin
        btb_5_pc <= btb_15_pc;
      end else if (4'he == io_aw_addr) begin
        btb_5_pc <= btb_14_pc;
      end else begin
        btb_5_pc <= _GEN_406;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_5_inst <= 32'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_5_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin
        btb_5_inst <= btb_15_inst;
      end else if (4'he == io_aw_addr) begin
        btb_5_inst <= btb_14_inst;
      end else begin
        btb_5_inst <= _GEN_407;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_5_exception_type <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_5_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin
        btb_5_exception_type <= btb_15_exception_type;
      end else if (4'he == io_aw_addr) begin
        btb_5_exception_type <= btb_14_exception_type;
      end else begin
        btb_5_exception_type <= _GEN_408;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_5_pre_pc_target <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_5_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin
        btb_5_pre_pc_target <= btb_15_pre_pc_target;
      end else if (4'he == io_aw_addr) begin
        btb_5_pre_pc_target <= btb_14_pre_pc_target;
      end else begin
        btb_5_pre_pc_target <= _GEN_409;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_5_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_5_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin
        btb_5_pre_lookup_data <= btb_15_pre_lookup_data;
      end else if (4'he == io_aw_addr) begin
        btb_5_pre_lookup_data <= btb_14_pre_lookup_data;
      end else begin
        btb_5_pre_lookup_data <= _GEN_410;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_5_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_5_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin
        btb_5_pre_hashcode <= btb_15_pre_hashcode;
      end else if (4'he == io_aw_addr) begin
        btb_5_pre_hashcode <= btb_14_pre_hashcode;
      end else begin
        btb_5_pre_hashcode <= _GEN_411;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_5_pre_pht <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_5_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin
        btb_5_pre_pht <= btb_15_pre_pht;
      end else if (4'he == io_aw_addr) begin
        btb_5_pre_pht <= btb_14_pre_pht;
      end else begin
        btb_5_pre_pht <= _GEN_412;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_5_pre_bht <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_5_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin
        btb_5_pre_bht <= btb_15_pre_bht;
      end else if (4'he == io_aw_addr) begin
        btb_5_pre_bht <= btb_14_pre_bht;
      end else begin
        btb_5_pre_bht <= _GEN_413;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_5_pre_lookup_value <= 8'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_5_pre_lookup_value <= io_in_pre_lookup_value;
      end else if (4'hf == io_aw_addr) begin
        btb_5_pre_lookup_value <= btb_15_pre_lookup_value;
      end else if (4'he == io_aw_addr) begin
        btb_5_pre_lookup_value <= btb_14_pre_lookup_value;
      end else begin
        btb_5_pre_lookup_value <= _GEN_414;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_5_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_5_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin
        btb_5_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag;
      end else if (4'he == io_aw_addr) begin
        btb_5_pre_decoder_branchD_flag <= btb_14_pre_decoder_branchD_flag;
      end else begin
        btb_5_pre_decoder_branchD_flag <= _GEN_415;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_5_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_5_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin
        btb_5_pre_decoder_jump <= btb_15_pre_decoder_jump;
      end else if (4'he == io_aw_addr) begin
        btb_5_pre_decoder_jump <= btb_14_pre_decoder_jump;
      end else begin
        btb_5_pre_decoder_jump <= _GEN_416;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_5_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_5_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin
        btb_5_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata;
      end else if (4'he == io_aw_addr) begin
        btb_5_pre_decoder_branchdata <= btb_14_pre_decoder_branchdata;
      end else begin
        btb_5_pre_decoder_branchdata <= _GEN_417;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_5_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_5_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin
        btb_5_pre_decoder_jr <= btb_15_pre_decoder_jr;
      end else if (4'he == io_aw_addr) begin
        btb_5_pre_decoder_jr <= btb_14_pre_decoder_jr;
      end else begin
        btb_5_pre_decoder_jr <= _GEN_418;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_5_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_5_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin
        btb_5_true_branch_state <= btb_15_true_branch_state;
      end else if (4'he == io_aw_addr) begin
        btb_5_true_branch_state <= btb_14_true_branch_state;
      end else begin
        btb_5_true_branch_state <= _GEN_419;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_6_pc <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_6_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin
        btb_6_pc <= btb_15_pc;
      end else if (4'he == io_aw_addr) begin
        btb_6_pc <= btb_14_pc;
      end else begin
        btb_6_pc <= _GEN_406;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_6_inst <= 32'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_6_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin
        btb_6_inst <= btb_15_inst;
      end else if (4'he == io_aw_addr) begin
        btb_6_inst <= btb_14_inst;
      end else begin
        btb_6_inst <= _GEN_407;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_6_exception_type <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_6_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin
        btb_6_exception_type <= btb_15_exception_type;
      end else if (4'he == io_aw_addr) begin
        btb_6_exception_type <= btb_14_exception_type;
      end else begin
        btb_6_exception_type <= _GEN_408;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_6_pre_pc_target <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_6_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin
        btb_6_pre_pc_target <= btb_15_pre_pc_target;
      end else if (4'he == io_aw_addr) begin
        btb_6_pre_pc_target <= btb_14_pre_pc_target;
      end else begin
        btb_6_pre_pc_target <= _GEN_409;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_6_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_6_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin
        btb_6_pre_lookup_data <= btb_15_pre_lookup_data;
      end else if (4'he == io_aw_addr) begin
        btb_6_pre_lookup_data <= btb_14_pre_lookup_data;
      end else begin
        btb_6_pre_lookup_data <= _GEN_410;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_6_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_6_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin
        btb_6_pre_hashcode <= btb_15_pre_hashcode;
      end else if (4'he == io_aw_addr) begin
        btb_6_pre_hashcode <= btb_14_pre_hashcode;
      end else begin
        btb_6_pre_hashcode <= _GEN_411;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_6_pre_pht <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_6_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin
        btb_6_pre_pht <= btb_15_pre_pht;
      end else if (4'he == io_aw_addr) begin
        btb_6_pre_pht <= btb_14_pre_pht;
      end else begin
        btb_6_pre_pht <= _GEN_412;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_6_pre_bht <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_6_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin
        btb_6_pre_bht <= btb_15_pre_bht;
      end else if (4'he == io_aw_addr) begin
        btb_6_pre_bht <= btb_14_pre_bht;
      end else begin
        btb_6_pre_bht <= _GEN_413;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_6_pre_lookup_value <= 8'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_6_pre_lookup_value <= io_in_pre_lookup_value;
      end else if (4'hf == io_aw_addr) begin
        btb_6_pre_lookup_value <= btb_15_pre_lookup_value;
      end else if (4'he == io_aw_addr) begin
        btb_6_pre_lookup_value <= btb_14_pre_lookup_value;
      end else begin
        btb_6_pre_lookup_value <= _GEN_414;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_6_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_6_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin
        btb_6_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag;
      end else if (4'he == io_aw_addr) begin
        btb_6_pre_decoder_branchD_flag <= btb_14_pre_decoder_branchD_flag;
      end else begin
        btb_6_pre_decoder_branchD_flag <= _GEN_415;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_6_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_6_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin
        btb_6_pre_decoder_jump <= btb_15_pre_decoder_jump;
      end else if (4'he == io_aw_addr) begin
        btb_6_pre_decoder_jump <= btb_14_pre_decoder_jump;
      end else begin
        btb_6_pre_decoder_jump <= _GEN_416;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_6_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_6_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin
        btb_6_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata;
      end else if (4'he == io_aw_addr) begin
        btb_6_pre_decoder_branchdata <= btb_14_pre_decoder_branchdata;
      end else begin
        btb_6_pre_decoder_branchdata <= _GEN_417;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_6_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_6_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin
        btb_6_pre_decoder_jr <= btb_15_pre_decoder_jr;
      end else if (4'he == io_aw_addr) begin
        btb_6_pre_decoder_jr <= btb_14_pre_decoder_jr;
      end else begin
        btb_6_pre_decoder_jr <= _GEN_418;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_6_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_6_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin
        btb_6_true_branch_state <= btb_15_true_branch_state;
      end else if (4'he == io_aw_addr) begin
        btb_6_true_branch_state <= btb_14_true_branch_state;
      end else begin
        btb_6_true_branch_state <= _GEN_419;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_7_pc <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_7_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin
        btb_7_pc <= btb_15_pc;
      end else if (4'he == io_aw_addr) begin
        btb_7_pc <= btb_14_pc;
      end else begin
        btb_7_pc <= _GEN_406;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_7_inst <= 32'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_7_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin
        btb_7_inst <= btb_15_inst;
      end else if (4'he == io_aw_addr) begin
        btb_7_inst <= btb_14_inst;
      end else begin
        btb_7_inst <= _GEN_407;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_7_exception_type <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_7_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin
        btb_7_exception_type <= btb_15_exception_type;
      end else if (4'he == io_aw_addr) begin
        btb_7_exception_type <= btb_14_exception_type;
      end else begin
        btb_7_exception_type <= _GEN_408;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_7_pre_pc_target <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_7_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin
        btb_7_pre_pc_target <= btb_15_pre_pc_target;
      end else if (4'he == io_aw_addr) begin
        btb_7_pre_pc_target <= btb_14_pre_pc_target;
      end else begin
        btb_7_pre_pc_target <= _GEN_409;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_7_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_7_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin
        btb_7_pre_lookup_data <= btb_15_pre_lookup_data;
      end else if (4'he == io_aw_addr) begin
        btb_7_pre_lookup_data <= btb_14_pre_lookup_data;
      end else begin
        btb_7_pre_lookup_data <= _GEN_410;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_7_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_7_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin
        btb_7_pre_hashcode <= btb_15_pre_hashcode;
      end else if (4'he == io_aw_addr) begin
        btb_7_pre_hashcode <= btb_14_pre_hashcode;
      end else begin
        btb_7_pre_hashcode <= _GEN_411;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_7_pre_pht <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_7_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin
        btb_7_pre_pht <= btb_15_pre_pht;
      end else if (4'he == io_aw_addr) begin
        btb_7_pre_pht <= btb_14_pre_pht;
      end else begin
        btb_7_pre_pht <= _GEN_412;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_7_pre_bht <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_7_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin
        btb_7_pre_bht <= btb_15_pre_bht;
      end else if (4'he == io_aw_addr) begin
        btb_7_pre_bht <= btb_14_pre_bht;
      end else begin
        btb_7_pre_bht <= _GEN_413;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_7_pre_lookup_value <= 8'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_7_pre_lookup_value <= io_in_pre_lookup_value;
      end else if (4'hf == io_aw_addr) begin
        btb_7_pre_lookup_value <= btb_15_pre_lookup_value;
      end else if (4'he == io_aw_addr) begin
        btb_7_pre_lookup_value <= btb_14_pre_lookup_value;
      end else begin
        btb_7_pre_lookup_value <= _GEN_414;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_7_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_7_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin
        btb_7_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag;
      end else if (4'he == io_aw_addr) begin
        btb_7_pre_decoder_branchD_flag <= btb_14_pre_decoder_branchD_flag;
      end else begin
        btb_7_pre_decoder_branchD_flag <= _GEN_415;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_7_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_7_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin
        btb_7_pre_decoder_jump <= btb_15_pre_decoder_jump;
      end else if (4'he == io_aw_addr) begin
        btb_7_pre_decoder_jump <= btb_14_pre_decoder_jump;
      end else begin
        btb_7_pre_decoder_jump <= _GEN_416;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_7_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_7_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin
        btb_7_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata;
      end else if (4'he == io_aw_addr) begin
        btb_7_pre_decoder_branchdata <= btb_14_pre_decoder_branchdata;
      end else begin
        btb_7_pre_decoder_branchdata <= _GEN_417;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_7_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_7_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin
        btb_7_pre_decoder_jr <= btb_15_pre_decoder_jr;
      end else if (4'he == io_aw_addr) begin
        btb_7_pre_decoder_jr <= btb_14_pre_decoder_jr;
      end else begin
        btb_7_pre_decoder_jr <= _GEN_418;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_7_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_7_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin
        btb_7_true_branch_state <= btb_15_true_branch_state;
      end else if (4'he == io_aw_addr) begin
        btb_7_true_branch_state <= btb_14_true_branch_state;
      end else begin
        btb_7_true_branch_state <= _GEN_419;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_8_pc <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_8_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin
        btb_8_pc <= btb_15_pc;
      end else if (4'he == io_aw_addr) begin
        btb_8_pc <= btb_14_pc;
      end else begin
        btb_8_pc <= _GEN_406;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_8_inst <= 32'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_8_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin
        btb_8_inst <= btb_15_inst;
      end else if (4'he == io_aw_addr) begin
        btb_8_inst <= btb_14_inst;
      end else begin
        btb_8_inst <= _GEN_407;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_8_exception_type <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_8_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin
        btb_8_exception_type <= btb_15_exception_type;
      end else if (4'he == io_aw_addr) begin
        btb_8_exception_type <= btb_14_exception_type;
      end else begin
        btb_8_exception_type <= _GEN_408;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_8_pre_pc_target <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_8_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin
        btb_8_pre_pc_target <= btb_15_pre_pc_target;
      end else if (4'he == io_aw_addr) begin
        btb_8_pre_pc_target <= btb_14_pre_pc_target;
      end else begin
        btb_8_pre_pc_target <= _GEN_409;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_8_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_8_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin
        btb_8_pre_lookup_data <= btb_15_pre_lookup_data;
      end else if (4'he == io_aw_addr) begin
        btb_8_pre_lookup_data <= btb_14_pre_lookup_data;
      end else begin
        btb_8_pre_lookup_data <= _GEN_410;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_8_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_8_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin
        btb_8_pre_hashcode <= btb_15_pre_hashcode;
      end else if (4'he == io_aw_addr) begin
        btb_8_pre_hashcode <= btb_14_pre_hashcode;
      end else begin
        btb_8_pre_hashcode <= _GEN_411;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_8_pre_pht <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_8_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin
        btb_8_pre_pht <= btb_15_pre_pht;
      end else if (4'he == io_aw_addr) begin
        btb_8_pre_pht <= btb_14_pre_pht;
      end else begin
        btb_8_pre_pht <= _GEN_412;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_8_pre_bht <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_8_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin
        btb_8_pre_bht <= btb_15_pre_bht;
      end else if (4'he == io_aw_addr) begin
        btb_8_pre_bht <= btb_14_pre_bht;
      end else begin
        btb_8_pre_bht <= _GEN_413;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_8_pre_lookup_value <= 8'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_8_pre_lookup_value <= io_in_pre_lookup_value;
      end else if (4'hf == io_aw_addr) begin
        btb_8_pre_lookup_value <= btb_15_pre_lookup_value;
      end else if (4'he == io_aw_addr) begin
        btb_8_pre_lookup_value <= btb_14_pre_lookup_value;
      end else begin
        btb_8_pre_lookup_value <= _GEN_414;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_8_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_8_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin
        btb_8_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag;
      end else if (4'he == io_aw_addr) begin
        btb_8_pre_decoder_branchD_flag <= btb_14_pre_decoder_branchD_flag;
      end else begin
        btb_8_pre_decoder_branchD_flag <= _GEN_415;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_8_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_8_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin
        btb_8_pre_decoder_jump <= btb_15_pre_decoder_jump;
      end else if (4'he == io_aw_addr) begin
        btb_8_pre_decoder_jump <= btb_14_pre_decoder_jump;
      end else begin
        btb_8_pre_decoder_jump <= _GEN_416;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_8_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_8_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin
        btb_8_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata;
      end else if (4'he == io_aw_addr) begin
        btb_8_pre_decoder_branchdata <= btb_14_pre_decoder_branchdata;
      end else begin
        btb_8_pre_decoder_branchdata <= _GEN_417;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_8_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_8_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin
        btb_8_pre_decoder_jr <= btb_15_pre_decoder_jr;
      end else if (4'he == io_aw_addr) begin
        btb_8_pre_decoder_jr <= btb_14_pre_decoder_jr;
      end else begin
        btb_8_pre_decoder_jr <= _GEN_418;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_8_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_8_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin
        btb_8_true_branch_state <= btb_15_true_branch_state;
      end else if (4'he == io_aw_addr) begin
        btb_8_true_branch_state <= btb_14_true_branch_state;
      end else begin
        btb_8_true_branch_state <= _GEN_419;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_9_pc <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_9_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin
        btb_9_pc <= btb_15_pc;
      end else if (4'he == io_aw_addr) begin
        btb_9_pc <= btb_14_pc;
      end else begin
        btb_9_pc <= _GEN_406;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_9_inst <= 32'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_9_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin
        btb_9_inst <= btb_15_inst;
      end else if (4'he == io_aw_addr) begin
        btb_9_inst <= btb_14_inst;
      end else begin
        btb_9_inst <= _GEN_407;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_9_exception_type <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_9_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin
        btb_9_exception_type <= btb_15_exception_type;
      end else if (4'he == io_aw_addr) begin
        btb_9_exception_type <= btb_14_exception_type;
      end else begin
        btb_9_exception_type <= _GEN_408;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_9_pre_pc_target <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_9_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin
        btb_9_pre_pc_target <= btb_15_pre_pc_target;
      end else if (4'he == io_aw_addr) begin
        btb_9_pre_pc_target <= btb_14_pre_pc_target;
      end else begin
        btb_9_pre_pc_target <= _GEN_409;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_9_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_9_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin
        btb_9_pre_lookup_data <= btb_15_pre_lookup_data;
      end else if (4'he == io_aw_addr) begin
        btb_9_pre_lookup_data <= btb_14_pre_lookup_data;
      end else begin
        btb_9_pre_lookup_data <= _GEN_410;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_9_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_9_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin
        btb_9_pre_hashcode <= btb_15_pre_hashcode;
      end else if (4'he == io_aw_addr) begin
        btb_9_pre_hashcode <= btb_14_pre_hashcode;
      end else begin
        btb_9_pre_hashcode <= _GEN_411;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_9_pre_pht <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_9_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin
        btb_9_pre_pht <= btb_15_pre_pht;
      end else if (4'he == io_aw_addr) begin
        btb_9_pre_pht <= btb_14_pre_pht;
      end else begin
        btb_9_pre_pht <= _GEN_412;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_9_pre_bht <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_9_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin
        btb_9_pre_bht <= btb_15_pre_bht;
      end else if (4'he == io_aw_addr) begin
        btb_9_pre_bht <= btb_14_pre_bht;
      end else begin
        btb_9_pre_bht <= _GEN_413;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_9_pre_lookup_value <= 8'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_9_pre_lookup_value <= io_in_pre_lookup_value;
      end else if (4'hf == io_aw_addr) begin
        btb_9_pre_lookup_value <= btb_15_pre_lookup_value;
      end else if (4'he == io_aw_addr) begin
        btb_9_pre_lookup_value <= btb_14_pre_lookup_value;
      end else begin
        btb_9_pre_lookup_value <= _GEN_414;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_9_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_9_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin
        btb_9_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag;
      end else if (4'he == io_aw_addr) begin
        btb_9_pre_decoder_branchD_flag <= btb_14_pre_decoder_branchD_flag;
      end else begin
        btb_9_pre_decoder_branchD_flag <= _GEN_415;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_9_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_9_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin
        btb_9_pre_decoder_jump <= btb_15_pre_decoder_jump;
      end else if (4'he == io_aw_addr) begin
        btb_9_pre_decoder_jump <= btb_14_pre_decoder_jump;
      end else begin
        btb_9_pre_decoder_jump <= _GEN_416;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_9_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_9_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin
        btb_9_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata;
      end else if (4'he == io_aw_addr) begin
        btb_9_pre_decoder_branchdata <= btb_14_pre_decoder_branchdata;
      end else begin
        btb_9_pre_decoder_branchdata <= _GEN_417;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_9_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_9_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin
        btb_9_pre_decoder_jr <= btb_15_pre_decoder_jr;
      end else if (4'he == io_aw_addr) begin
        btb_9_pre_decoder_jr <= btb_14_pre_decoder_jr;
      end else begin
        btb_9_pre_decoder_jr <= _GEN_418;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_9_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_9_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin
        btb_9_true_branch_state <= btb_15_true_branch_state;
      end else if (4'he == io_aw_addr) begin
        btb_9_true_branch_state <= btb_14_true_branch_state;
      end else begin
        btb_9_true_branch_state <= _GEN_419;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_10_pc <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_10_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin
        btb_10_pc <= btb_15_pc;
      end else if (4'he == io_aw_addr) begin
        btb_10_pc <= btb_14_pc;
      end else begin
        btb_10_pc <= _GEN_406;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_10_inst <= 32'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_10_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin
        btb_10_inst <= btb_15_inst;
      end else if (4'he == io_aw_addr) begin
        btb_10_inst <= btb_14_inst;
      end else begin
        btb_10_inst <= _GEN_407;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_10_exception_type <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_10_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin
        btb_10_exception_type <= btb_15_exception_type;
      end else if (4'he == io_aw_addr) begin
        btb_10_exception_type <= btb_14_exception_type;
      end else begin
        btb_10_exception_type <= _GEN_408;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_10_pre_pc_target <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_10_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin
        btb_10_pre_pc_target <= btb_15_pre_pc_target;
      end else if (4'he == io_aw_addr) begin
        btb_10_pre_pc_target <= btb_14_pre_pc_target;
      end else begin
        btb_10_pre_pc_target <= _GEN_409;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_10_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_10_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin
        btb_10_pre_lookup_data <= btb_15_pre_lookup_data;
      end else if (4'he == io_aw_addr) begin
        btb_10_pre_lookup_data <= btb_14_pre_lookup_data;
      end else begin
        btb_10_pre_lookup_data <= _GEN_410;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_10_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_10_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin
        btb_10_pre_hashcode <= btb_15_pre_hashcode;
      end else if (4'he == io_aw_addr) begin
        btb_10_pre_hashcode <= btb_14_pre_hashcode;
      end else begin
        btb_10_pre_hashcode <= _GEN_411;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_10_pre_pht <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_10_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin
        btb_10_pre_pht <= btb_15_pre_pht;
      end else if (4'he == io_aw_addr) begin
        btb_10_pre_pht <= btb_14_pre_pht;
      end else begin
        btb_10_pre_pht <= _GEN_412;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_10_pre_bht <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_10_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin
        btb_10_pre_bht <= btb_15_pre_bht;
      end else if (4'he == io_aw_addr) begin
        btb_10_pre_bht <= btb_14_pre_bht;
      end else begin
        btb_10_pre_bht <= _GEN_413;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_10_pre_lookup_value <= 8'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_10_pre_lookup_value <= io_in_pre_lookup_value;
      end else if (4'hf == io_aw_addr) begin
        btb_10_pre_lookup_value <= btb_15_pre_lookup_value;
      end else if (4'he == io_aw_addr) begin
        btb_10_pre_lookup_value <= btb_14_pre_lookup_value;
      end else begin
        btb_10_pre_lookup_value <= _GEN_414;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_10_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_10_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin
        btb_10_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag;
      end else if (4'he == io_aw_addr) begin
        btb_10_pre_decoder_branchD_flag <= btb_14_pre_decoder_branchD_flag;
      end else begin
        btb_10_pre_decoder_branchD_flag <= _GEN_415;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_10_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_10_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin
        btb_10_pre_decoder_jump <= btb_15_pre_decoder_jump;
      end else if (4'he == io_aw_addr) begin
        btb_10_pre_decoder_jump <= btb_14_pre_decoder_jump;
      end else begin
        btb_10_pre_decoder_jump <= _GEN_416;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_10_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_10_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin
        btb_10_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata;
      end else if (4'he == io_aw_addr) begin
        btb_10_pre_decoder_branchdata <= btb_14_pre_decoder_branchdata;
      end else begin
        btb_10_pre_decoder_branchdata <= _GEN_417;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_10_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_10_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin
        btb_10_pre_decoder_jr <= btb_15_pre_decoder_jr;
      end else if (4'he == io_aw_addr) begin
        btb_10_pre_decoder_jr <= btb_14_pre_decoder_jr;
      end else begin
        btb_10_pre_decoder_jr <= _GEN_418;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_10_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'ha == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_10_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin
        btb_10_true_branch_state <= btb_15_true_branch_state;
      end else if (4'he == io_aw_addr) begin
        btb_10_true_branch_state <= btb_14_true_branch_state;
      end else begin
        btb_10_true_branch_state <= _GEN_419;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_11_pc <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_11_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin
        btb_11_pc <= btb_15_pc;
      end else if (4'he == io_aw_addr) begin
        btb_11_pc <= btb_14_pc;
      end else begin
        btb_11_pc <= _GEN_406;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_11_inst <= 32'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_11_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin
        btb_11_inst <= btb_15_inst;
      end else if (4'he == io_aw_addr) begin
        btb_11_inst <= btb_14_inst;
      end else begin
        btb_11_inst <= _GEN_407;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_11_exception_type <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_11_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin
        btb_11_exception_type <= btb_15_exception_type;
      end else if (4'he == io_aw_addr) begin
        btb_11_exception_type <= btb_14_exception_type;
      end else begin
        btb_11_exception_type <= _GEN_408;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_11_pre_pc_target <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_11_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin
        btb_11_pre_pc_target <= btb_15_pre_pc_target;
      end else if (4'he == io_aw_addr) begin
        btb_11_pre_pc_target <= btb_14_pre_pc_target;
      end else begin
        btb_11_pre_pc_target <= _GEN_409;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_11_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_11_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin
        btb_11_pre_lookup_data <= btb_15_pre_lookup_data;
      end else if (4'he == io_aw_addr) begin
        btb_11_pre_lookup_data <= btb_14_pre_lookup_data;
      end else begin
        btb_11_pre_lookup_data <= _GEN_410;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_11_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_11_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin
        btb_11_pre_hashcode <= btb_15_pre_hashcode;
      end else if (4'he == io_aw_addr) begin
        btb_11_pre_hashcode <= btb_14_pre_hashcode;
      end else begin
        btb_11_pre_hashcode <= _GEN_411;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_11_pre_pht <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_11_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin
        btb_11_pre_pht <= btb_15_pre_pht;
      end else if (4'he == io_aw_addr) begin
        btb_11_pre_pht <= btb_14_pre_pht;
      end else begin
        btb_11_pre_pht <= _GEN_412;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_11_pre_bht <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_11_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin
        btb_11_pre_bht <= btb_15_pre_bht;
      end else if (4'he == io_aw_addr) begin
        btb_11_pre_bht <= btb_14_pre_bht;
      end else begin
        btb_11_pre_bht <= _GEN_413;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_11_pre_lookup_value <= 8'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_11_pre_lookup_value <= io_in_pre_lookup_value;
      end else if (4'hf == io_aw_addr) begin
        btb_11_pre_lookup_value <= btb_15_pre_lookup_value;
      end else if (4'he == io_aw_addr) begin
        btb_11_pre_lookup_value <= btb_14_pre_lookup_value;
      end else begin
        btb_11_pre_lookup_value <= _GEN_414;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_11_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_11_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin
        btb_11_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag;
      end else if (4'he == io_aw_addr) begin
        btb_11_pre_decoder_branchD_flag <= btb_14_pre_decoder_branchD_flag;
      end else begin
        btb_11_pre_decoder_branchD_flag <= _GEN_415;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_11_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_11_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin
        btb_11_pre_decoder_jump <= btb_15_pre_decoder_jump;
      end else if (4'he == io_aw_addr) begin
        btb_11_pre_decoder_jump <= btb_14_pre_decoder_jump;
      end else begin
        btb_11_pre_decoder_jump <= _GEN_416;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_11_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_11_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin
        btb_11_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata;
      end else if (4'he == io_aw_addr) begin
        btb_11_pre_decoder_branchdata <= btb_14_pre_decoder_branchdata;
      end else begin
        btb_11_pre_decoder_branchdata <= _GEN_417;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_11_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_11_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin
        btb_11_pre_decoder_jr <= btb_15_pre_decoder_jr;
      end else if (4'he == io_aw_addr) begin
        btb_11_pre_decoder_jr <= btb_14_pre_decoder_jr;
      end else begin
        btb_11_pre_decoder_jr <= _GEN_418;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_11_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hb == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_11_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin
        btb_11_true_branch_state <= btb_15_true_branch_state;
      end else if (4'he == io_aw_addr) begin
        btb_11_true_branch_state <= btb_14_true_branch_state;
      end else begin
        btb_11_true_branch_state <= _GEN_419;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_12_pc <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_12_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin
        btb_12_pc <= btb_15_pc;
      end else if (4'he == io_aw_addr) begin
        btb_12_pc <= btb_14_pc;
      end else begin
        btb_12_pc <= _GEN_406;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_12_inst <= 32'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_12_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin
        btb_12_inst <= btb_15_inst;
      end else if (4'he == io_aw_addr) begin
        btb_12_inst <= btb_14_inst;
      end else begin
        btb_12_inst <= _GEN_407;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_12_exception_type <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_12_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin
        btb_12_exception_type <= btb_15_exception_type;
      end else if (4'he == io_aw_addr) begin
        btb_12_exception_type <= btb_14_exception_type;
      end else begin
        btb_12_exception_type <= _GEN_408;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_12_pre_pc_target <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_12_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin
        btb_12_pre_pc_target <= btb_15_pre_pc_target;
      end else if (4'he == io_aw_addr) begin
        btb_12_pre_pc_target <= btb_14_pre_pc_target;
      end else begin
        btb_12_pre_pc_target <= _GEN_409;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_12_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_12_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin
        btb_12_pre_lookup_data <= btb_15_pre_lookup_data;
      end else if (4'he == io_aw_addr) begin
        btb_12_pre_lookup_data <= btb_14_pre_lookup_data;
      end else begin
        btb_12_pre_lookup_data <= _GEN_410;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_12_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_12_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin
        btb_12_pre_hashcode <= btb_15_pre_hashcode;
      end else if (4'he == io_aw_addr) begin
        btb_12_pre_hashcode <= btb_14_pre_hashcode;
      end else begin
        btb_12_pre_hashcode <= _GEN_411;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_12_pre_pht <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_12_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin
        btb_12_pre_pht <= btb_15_pre_pht;
      end else if (4'he == io_aw_addr) begin
        btb_12_pre_pht <= btb_14_pre_pht;
      end else begin
        btb_12_pre_pht <= _GEN_412;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_12_pre_bht <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_12_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin
        btb_12_pre_bht <= btb_15_pre_bht;
      end else if (4'he == io_aw_addr) begin
        btb_12_pre_bht <= btb_14_pre_bht;
      end else begin
        btb_12_pre_bht <= _GEN_413;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_12_pre_lookup_value <= 8'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_12_pre_lookup_value <= io_in_pre_lookup_value;
      end else if (4'hf == io_aw_addr) begin
        btb_12_pre_lookup_value <= btb_15_pre_lookup_value;
      end else if (4'he == io_aw_addr) begin
        btb_12_pre_lookup_value <= btb_14_pre_lookup_value;
      end else begin
        btb_12_pre_lookup_value <= _GEN_414;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_12_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_12_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin
        btb_12_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag;
      end else if (4'he == io_aw_addr) begin
        btb_12_pre_decoder_branchD_flag <= btb_14_pre_decoder_branchD_flag;
      end else begin
        btb_12_pre_decoder_branchD_flag <= _GEN_415;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_12_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_12_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin
        btb_12_pre_decoder_jump <= btb_15_pre_decoder_jump;
      end else if (4'he == io_aw_addr) begin
        btb_12_pre_decoder_jump <= btb_14_pre_decoder_jump;
      end else begin
        btb_12_pre_decoder_jump <= _GEN_416;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_12_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_12_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin
        btb_12_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata;
      end else if (4'he == io_aw_addr) begin
        btb_12_pre_decoder_branchdata <= btb_14_pre_decoder_branchdata;
      end else begin
        btb_12_pre_decoder_branchdata <= _GEN_417;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_12_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_12_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin
        btb_12_pre_decoder_jr <= btb_15_pre_decoder_jr;
      end else if (4'he == io_aw_addr) begin
        btb_12_pre_decoder_jr <= btb_14_pre_decoder_jr;
      end else begin
        btb_12_pre_decoder_jr <= _GEN_418;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_12_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hc == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_12_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin
        btb_12_true_branch_state <= btb_15_true_branch_state;
      end else if (4'he == io_aw_addr) begin
        btb_12_true_branch_state <= btb_14_true_branch_state;
      end else begin
        btb_12_true_branch_state <= _GEN_419;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_13_pc <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_13_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin
        btb_13_pc <= btb_15_pc;
      end else if (4'he == io_aw_addr) begin
        btb_13_pc <= btb_14_pc;
      end else begin
        btb_13_pc <= _GEN_406;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_13_inst <= 32'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_13_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin
        btb_13_inst <= btb_15_inst;
      end else if (4'he == io_aw_addr) begin
        btb_13_inst <= btb_14_inst;
      end else begin
        btb_13_inst <= _GEN_407;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_13_exception_type <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_13_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin
        btb_13_exception_type <= btb_15_exception_type;
      end else if (4'he == io_aw_addr) begin
        btb_13_exception_type <= btb_14_exception_type;
      end else begin
        btb_13_exception_type <= _GEN_408;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_13_pre_pc_target <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_13_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin
        btb_13_pre_pc_target <= btb_15_pre_pc_target;
      end else if (4'he == io_aw_addr) begin
        btb_13_pre_pc_target <= btb_14_pre_pc_target;
      end else begin
        btb_13_pre_pc_target <= _GEN_409;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_13_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_13_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin
        btb_13_pre_lookup_data <= btb_15_pre_lookup_data;
      end else if (4'he == io_aw_addr) begin
        btb_13_pre_lookup_data <= btb_14_pre_lookup_data;
      end else begin
        btb_13_pre_lookup_data <= _GEN_410;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_13_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_13_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin
        btb_13_pre_hashcode <= btb_15_pre_hashcode;
      end else if (4'he == io_aw_addr) begin
        btb_13_pre_hashcode <= btb_14_pre_hashcode;
      end else begin
        btb_13_pre_hashcode <= _GEN_411;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_13_pre_pht <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_13_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin
        btb_13_pre_pht <= btb_15_pre_pht;
      end else if (4'he == io_aw_addr) begin
        btb_13_pre_pht <= btb_14_pre_pht;
      end else begin
        btb_13_pre_pht <= _GEN_412;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_13_pre_bht <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_13_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin
        btb_13_pre_bht <= btb_15_pre_bht;
      end else if (4'he == io_aw_addr) begin
        btb_13_pre_bht <= btb_14_pre_bht;
      end else begin
        btb_13_pre_bht <= _GEN_413;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_13_pre_lookup_value <= 8'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_13_pre_lookup_value <= io_in_pre_lookup_value;
      end else if (4'hf == io_aw_addr) begin
        btb_13_pre_lookup_value <= btb_15_pre_lookup_value;
      end else if (4'he == io_aw_addr) begin
        btb_13_pre_lookup_value <= btb_14_pre_lookup_value;
      end else begin
        btb_13_pre_lookup_value <= _GEN_414;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_13_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_13_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin
        btb_13_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag;
      end else if (4'he == io_aw_addr) begin
        btb_13_pre_decoder_branchD_flag <= btb_14_pre_decoder_branchD_flag;
      end else begin
        btb_13_pre_decoder_branchD_flag <= _GEN_415;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_13_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_13_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin
        btb_13_pre_decoder_jump <= btb_15_pre_decoder_jump;
      end else if (4'he == io_aw_addr) begin
        btb_13_pre_decoder_jump <= btb_14_pre_decoder_jump;
      end else begin
        btb_13_pre_decoder_jump <= _GEN_416;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_13_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_13_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin
        btb_13_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata;
      end else if (4'he == io_aw_addr) begin
        btb_13_pre_decoder_branchdata <= btb_14_pre_decoder_branchdata;
      end else begin
        btb_13_pre_decoder_branchdata <= _GEN_417;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_13_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_13_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin
        btb_13_pre_decoder_jr <= btb_15_pre_decoder_jr;
      end else if (4'he == io_aw_addr) begin
        btb_13_pre_decoder_jr <= btb_14_pre_decoder_jr;
      end else begin
        btb_13_pre_decoder_jr <= _GEN_418;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_13_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hd == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_13_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin
        btb_13_true_branch_state <= btb_15_true_branch_state;
      end else if (4'he == io_aw_addr) begin
        btb_13_true_branch_state <= btb_14_true_branch_state;
      end else begin
        btb_13_true_branch_state <= _GEN_419;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_14_pc <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_14_pc <= io_in_pc;
      end else if (4'hf == io_aw_addr) begin
        btb_14_pc <= btb_15_pc;
      end else if (!(4'he == io_aw_addr)) begin
        btb_14_pc <= _GEN_406;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_14_inst <= 32'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_14_inst <= io_in_inst;
      end else if (4'hf == io_aw_addr) begin
        btb_14_inst <= btb_15_inst;
      end else if (!(4'he == io_aw_addr)) begin
        btb_14_inst <= _GEN_407;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_14_exception_type <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_14_exception_type <= 2'h0;
      end else if (4'hf == io_aw_addr) begin
        btb_14_exception_type <= btb_15_exception_type;
      end else if (!(4'he == io_aw_addr)) begin
        btb_14_exception_type <= _GEN_408;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_14_pre_pc_target <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_14_pre_pc_target <= io_in_pre_pc_target;
      end else if (4'hf == io_aw_addr) begin
        btb_14_pre_pc_target <= btb_15_pre_pc_target;
      end else if (!(4'he == io_aw_addr)) begin
        btb_14_pre_pc_target <= _GEN_409;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_14_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_14_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (4'hf == io_aw_addr) begin
        btb_14_pre_lookup_data <= btb_15_pre_lookup_data;
      end else if (!(4'he == io_aw_addr)) begin
        btb_14_pre_lookup_data <= _GEN_410;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_14_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_14_pre_hashcode <= io_in_pre_hashcode;
      end else if (4'hf == io_aw_addr) begin
        btb_14_pre_hashcode <= btb_15_pre_hashcode;
      end else if (!(4'he == io_aw_addr)) begin
        btb_14_pre_hashcode <= _GEN_411;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_14_pre_pht <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_14_pre_pht <= io_in_pre_pht;
      end else if (4'hf == io_aw_addr) begin
        btb_14_pre_pht <= btb_15_pre_pht;
      end else if (!(4'he == io_aw_addr)) begin
        btb_14_pre_pht <= _GEN_412;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_14_pre_bht <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_14_pre_bht <= io_in_pre_bht;
      end else if (4'hf == io_aw_addr) begin
        btb_14_pre_bht <= btb_15_pre_bht;
      end else if (!(4'he == io_aw_addr)) begin
        btb_14_pre_bht <= _GEN_413;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_14_pre_lookup_value <= 8'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_14_pre_lookup_value <= io_in_pre_lookup_value;
      end else if (4'hf == io_aw_addr) begin
        btb_14_pre_lookup_value <= btb_15_pre_lookup_value;
      end else if (!(4'he == io_aw_addr)) begin
        btb_14_pre_lookup_value <= _GEN_414;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_14_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_14_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (4'hf == io_aw_addr) begin
        btb_14_pre_decoder_branchD_flag <= btb_15_pre_decoder_branchD_flag;
      end else if (!(4'he == io_aw_addr)) begin
        btb_14_pre_decoder_branchD_flag <= _GEN_415;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_14_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_14_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (4'hf == io_aw_addr) begin
        btb_14_pre_decoder_jump <= btb_15_pre_decoder_jump;
      end else if (!(4'he == io_aw_addr)) begin
        btb_14_pre_decoder_jump <= _GEN_416;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_14_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_14_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (4'hf == io_aw_addr) begin
        btb_14_pre_decoder_branchdata <= btb_15_pre_decoder_branchdata;
      end else if (!(4'he == io_aw_addr)) begin
        btb_14_pre_decoder_branchdata <= _GEN_417;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_14_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_14_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (4'hf == io_aw_addr) begin
        btb_14_pre_decoder_jr <= btb_15_pre_decoder_jr;
      end else if (!(4'he == io_aw_addr)) begin
        btb_14_pre_decoder_jr <= _GEN_418;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_14_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'he == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_14_true_branch_state <= io_in_true_branch_state;
      end else if (4'hf == io_aw_addr) begin
        btb_14_true_branch_state <= btb_15_true_branch_state;
      end else if (!(4'he == io_aw_addr)) begin
        btb_14_true_branch_state <= _GEN_419;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_15_pc <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_15_pc <= io_in_pc;
      end else if (!(4'hf == io_aw_addr)) begin
        if (4'he == io_aw_addr) begin
          btb_15_pc <= btb_14_pc;
        end else begin
          btb_15_pc <= _GEN_406;
        end
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_15_inst <= 32'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_15_inst <= io_in_inst;
      end else if (!(4'hf == io_aw_addr)) begin
        if (4'he == io_aw_addr) begin
          btb_15_inst <= btb_14_inst;
        end else begin
          btb_15_inst <= _GEN_407;
        end
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_15_exception_type <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_15_exception_type <= 2'h0;
      end else if (!(4'hf == io_aw_addr)) begin
        if (4'he == io_aw_addr) begin
          btb_15_exception_type <= btb_14_exception_type;
        end else begin
          btb_15_exception_type <= _GEN_408;
        end
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_15_pre_pc_target <= 64'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_15_pre_pc_target <= io_in_pre_pc_target;
      end else if (!(4'hf == io_aw_addr)) begin
        if (4'he == io_aw_addr) begin
          btb_15_pre_pc_target <= btb_14_pre_pc_target;
        end else begin
          btb_15_pre_pc_target <= _GEN_409;
        end
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_15_pre_lookup_data <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_15_pre_lookup_data <= io_in_pre_lookup_data;
      end else if (!(4'hf == io_aw_addr)) begin
        if (4'he == io_aw_addr) begin
          btb_15_pre_lookup_data <= btb_14_pre_lookup_data;
        end else begin
          btb_15_pre_lookup_data <= _GEN_410;
        end
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_15_pre_hashcode <= 4'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_15_pre_hashcode <= io_in_pre_hashcode;
      end else if (!(4'hf == io_aw_addr)) begin
        if (4'he == io_aw_addr) begin
          btb_15_pre_hashcode <= btb_14_pre_hashcode;
        end else begin
          btb_15_pre_hashcode <= _GEN_411;
        end
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_15_pre_pht <= 2'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_15_pre_pht <= io_in_pre_pht;
      end else if (!(4'hf == io_aw_addr)) begin
        if (4'he == io_aw_addr) begin
          btb_15_pre_pht <= btb_14_pre_pht;
        end else begin
          btb_15_pre_pht <= _GEN_412;
        end
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_15_pre_bht <= 7'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_15_pre_bht <= io_in_pre_bht;
      end else if (!(4'hf == io_aw_addr)) begin
        if (4'he == io_aw_addr) begin
          btb_15_pre_bht <= btb_14_pre_bht;
        end else begin
          btb_15_pre_bht <= _GEN_413;
        end
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_15_pre_lookup_value <= 8'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_15_pre_lookup_value <= io_in_pre_lookup_value;
      end else if (!(4'hf == io_aw_addr)) begin
        if (4'he == io_aw_addr) begin
          btb_15_pre_lookup_value <= btb_14_pre_lookup_value;
        end else begin
          btb_15_pre_lookup_value <= _GEN_414;
        end
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_15_pre_decoder_branchD_flag <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_15_pre_decoder_branchD_flag <= io_in_pre_decoder_branchD_flag;
      end else if (!(4'hf == io_aw_addr)) begin
        if (4'he == io_aw_addr) begin
          btb_15_pre_decoder_branchD_flag <= btb_14_pre_decoder_branchD_flag;
        end else begin
          btb_15_pre_decoder_branchD_flag <= _GEN_415;
        end
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_15_pre_decoder_jump <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_15_pre_decoder_jump <= io_in_pre_decoder_jump;
      end else if (!(4'hf == io_aw_addr)) begin
        if (4'he == io_aw_addr) begin
          btb_15_pre_decoder_jump <= btb_14_pre_decoder_jump;
        end else begin
          btb_15_pre_decoder_jump <= _GEN_416;
        end
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_15_pre_decoder_branchdata <= 6'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_15_pre_decoder_branchdata <= io_in_pre_decoder_branchdata;
      end else if (!(4'hf == io_aw_addr)) begin
        if (4'he == io_aw_addr) begin
          btb_15_pre_decoder_branchdata <= btb_14_pre_decoder_branchdata;
        end else begin
          btb_15_pre_decoder_branchdata <= _GEN_417;
        end
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_15_pre_decoder_jr <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_15_pre_decoder_jr <= io_in_pre_decoder_jr;
      end else if (!(4'hf == io_aw_addr)) begin
        if (4'he == io_aw_addr) begin
          btb_15_pre_decoder_jr <= btb_14_pre_decoder_jr;
        end else begin
          btb_15_pre_decoder_jr <= _GEN_418;
        end
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 107:21]
      btb_15_true_branch_state <= 1'h0; // @[ports_lookup_table.scala 107:{27,27,27,27,27}]
    end else if (4'hf == io_aw_addr) begin // @[ports_lookup_table.scala 105:22]
      if (io_write) begin
        btb_15_true_branch_state <= io_in_true_branch_state;
      end else if (!(4'hf == io_aw_addr)) begin
        if (4'he == io_aw_addr) begin
          btb_15_true_branch_state <= btb_14_true_branch_state;
        end else begin
          btb_15_true_branch_state <= _GEN_419;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  btb_0_pc = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  btb_0_inst = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  btb_0_exception_type = _RAND_2[1:0];
  _RAND_3 = {2{`RANDOM}};
  btb_0_pre_pc_target = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  btb_0_pre_lookup_data = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  btb_0_pre_hashcode = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  btb_0_pre_pht = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  btb_0_pre_bht = _RAND_7[6:0];
  _RAND_8 = {1{`RANDOM}};
  btb_0_pre_lookup_value = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  btb_0_pre_decoder_branchD_flag = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  btb_0_pre_decoder_jump = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  btb_0_pre_decoder_branchdata = _RAND_11[5:0];
  _RAND_12 = {1{`RANDOM}};
  btb_0_pre_decoder_jr = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  btb_0_true_branch_state = _RAND_13[0:0];
  _RAND_14 = {2{`RANDOM}};
  btb_1_pc = _RAND_14[63:0];
  _RAND_15 = {1{`RANDOM}};
  btb_1_inst = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  btb_1_exception_type = _RAND_16[1:0];
  _RAND_17 = {2{`RANDOM}};
  btb_1_pre_pc_target = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  btb_1_pre_lookup_data = _RAND_18[6:0];
  _RAND_19 = {1{`RANDOM}};
  btb_1_pre_hashcode = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  btb_1_pre_pht = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  btb_1_pre_bht = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  btb_1_pre_lookup_value = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  btb_1_pre_decoder_branchD_flag = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  btb_1_pre_decoder_jump = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  btb_1_pre_decoder_branchdata = _RAND_25[5:0];
  _RAND_26 = {1{`RANDOM}};
  btb_1_pre_decoder_jr = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  btb_1_true_branch_state = _RAND_27[0:0];
  _RAND_28 = {2{`RANDOM}};
  btb_2_pc = _RAND_28[63:0];
  _RAND_29 = {1{`RANDOM}};
  btb_2_inst = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  btb_2_exception_type = _RAND_30[1:0];
  _RAND_31 = {2{`RANDOM}};
  btb_2_pre_pc_target = _RAND_31[63:0];
  _RAND_32 = {1{`RANDOM}};
  btb_2_pre_lookup_data = _RAND_32[6:0];
  _RAND_33 = {1{`RANDOM}};
  btb_2_pre_hashcode = _RAND_33[3:0];
  _RAND_34 = {1{`RANDOM}};
  btb_2_pre_pht = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  btb_2_pre_bht = _RAND_35[6:0];
  _RAND_36 = {1{`RANDOM}};
  btb_2_pre_lookup_value = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  btb_2_pre_decoder_branchD_flag = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  btb_2_pre_decoder_jump = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  btb_2_pre_decoder_branchdata = _RAND_39[5:0];
  _RAND_40 = {1{`RANDOM}};
  btb_2_pre_decoder_jr = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  btb_2_true_branch_state = _RAND_41[0:0];
  _RAND_42 = {2{`RANDOM}};
  btb_3_pc = _RAND_42[63:0];
  _RAND_43 = {1{`RANDOM}};
  btb_3_inst = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  btb_3_exception_type = _RAND_44[1:0];
  _RAND_45 = {2{`RANDOM}};
  btb_3_pre_pc_target = _RAND_45[63:0];
  _RAND_46 = {1{`RANDOM}};
  btb_3_pre_lookup_data = _RAND_46[6:0];
  _RAND_47 = {1{`RANDOM}};
  btb_3_pre_hashcode = _RAND_47[3:0];
  _RAND_48 = {1{`RANDOM}};
  btb_3_pre_pht = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  btb_3_pre_bht = _RAND_49[6:0];
  _RAND_50 = {1{`RANDOM}};
  btb_3_pre_lookup_value = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  btb_3_pre_decoder_branchD_flag = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  btb_3_pre_decoder_jump = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  btb_3_pre_decoder_branchdata = _RAND_53[5:0];
  _RAND_54 = {1{`RANDOM}};
  btb_3_pre_decoder_jr = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  btb_3_true_branch_state = _RAND_55[0:0];
  _RAND_56 = {2{`RANDOM}};
  btb_4_pc = _RAND_56[63:0];
  _RAND_57 = {1{`RANDOM}};
  btb_4_inst = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  btb_4_exception_type = _RAND_58[1:0];
  _RAND_59 = {2{`RANDOM}};
  btb_4_pre_pc_target = _RAND_59[63:0];
  _RAND_60 = {1{`RANDOM}};
  btb_4_pre_lookup_data = _RAND_60[6:0];
  _RAND_61 = {1{`RANDOM}};
  btb_4_pre_hashcode = _RAND_61[3:0];
  _RAND_62 = {1{`RANDOM}};
  btb_4_pre_pht = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  btb_4_pre_bht = _RAND_63[6:0];
  _RAND_64 = {1{`RANDOM}};
  btb_4_pre_lookup_value = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  btb_4_pre_decoder_branchD_flag = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  btb_4_pre_decoder_jump = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  btb_4_pre_decoder_branchdata = _RAND_67[5:0];
  _RAND_68 = {1{`RANDOM}};
  btb_4_pre_decoder_jr = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  btb_4_true_branch_state = _RAND_69[0:0];
  _RAND_70 = {2{`RANDOM}};
  btb_5_pc = _RAND_70[63:0];
  _RAND_71 = {1{`RANDOM}};
  btb_5_inst = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  btb_5_exception_type = _RAND_72[1:0];
  _RAND_73 = {2{`RANDOM}};
  btb_5_pre_pc_target = _RAND_73[63:0];
  _RAND_74 = {1{`RANDOM}};
  btb_5_pre_lookup_data = _RAND_74[6:0];
  _RAND_75 = {1{`RANDOM}};
  btb_5_pre_hashcode = _RAND_75[3:0];
  _RAND_76 = {1{`RANDOM}};
  btb_5_pre_pht = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  btb_5_pre_bht = _RAND_77[6:0];
  _RAND_78 = {1{`RANDOM}};
  btb_5_pre_lookup_value = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  btb_5_pre_decoder_branchD_flag = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  btb_5_pre_decoder_jump = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  btb_5_pre_decoder_branchdata = _RAND_81[5:0];
  _RAND_82 = {1{`RANDOM}};
  btb_5_pre_decoder_jr = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  btb_5_true_branch_state = _RAND_83[0:0];
  _RAND_84 = {2{`RANDOM}};
  btb_6_pc = _RAND_84[63:0];
  _RAND_85 = {1{`RANDOM}};
  btb_6_inst = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  btb_6_exception_type = _RAND_86[1:0];
  _RAND_87 = {2{`RANDOM}};
  btb_6_pre_pc_target = _RAND_87[63:0];
  _RAND_88 = {1{`RANDOM}};
  btb_6_pre_lookup_data = _RAND_88[6:0];
  _RAND_89 = {1{`RANDOM}};
  btb_6_pre_hashcode = _RAND_89[3:0];
  _RAND_90 = {1{`RANDOM}};
  btb_6_pre_pht = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  btb_6_pre_bht = _RAND_91[6:0];
  _RAND_92 = {1{`RANDOM}};
  btb_6_pre_lookup_value = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  btb_6_pre_decoder_branchD_flag = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  btb_6_pre_decoder_jump = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  btb_6_pre_decoder_branchdata = _RAND_95[5:0];
  _RAND_96 = {1{`RANDOM}};
  btb_6_pre_decoder_jr = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  btb_6_true_branch_state = _RAND_97[0:0];
  _RAND_98 = {2{`RANDOM}};
  btb_7_pc = _RAND_98[63:0];
  _RAND_99 = {1{`RANDOM}};
  btb_7_inst = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  btb_7_exception_type = _RAND_100[1:0];
  _RAND_101 = {2{`RANDOM}};
  btb_7_pre_pc_target = _RAND_101[63:0];
  _RAND_102 = {1{`RANDOM}};
  btb_7_pre_lookup_data = _RAND_102[6:0];
  _RAND_103 = {1{`RANDOM}};
  btb_7_pre_hashcode = _RAND_103[3:0];
  _RAND_104 = {1{`RANDOM}};
  btb_7_pre_pht = _RAND_104[1:0];
  _RAND_105 = {1{`RANDOM}};
  btb_7_pre_bht = _RAND_105[6:0];
  _RAND_106 = {1{`RANDOM}};
  btb_7_pre_lookup_value = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  btb_7_pre_decoder_branchD_flag = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  btb_7_pre_decoder_jump = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  btb_7_pre_decoder_branchdata = _RAND_109[5:0];
  _RAND_110 = {1{`RANDOM}};
  btb_7_pre_decoder_jr = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  btb_7_true_branch_state = _RAND_111[0:0];
  _RAND_112 = {2{`RANDOM}};
  btb_8_pc = _RAND_112[63:0];
  _RAND_113 = {1{`RANDOM}};
  btb_8_inst = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  btb_8_exception_type = _RAND_114[1:0];
  _RAND_115 = {2{`RANDOM}};
  btb_8_pre_pc_target = _RAND_115[63:0];
  _RAND_116 = {1{`RANDOM}};
  btb_8_pre_lookup_data = _RAND_116[6:0];
  _RAND_117 = {1{`RANDOM}};
  btb_8_pre_hashcode = _RAND_117[3:0];
  _RAND_118 = {1{`RANDOM}};
  btb_8_pre_pht = _RAND_118[1:0];
  _RAND_119 = {1{`RANDOM}};
  btb_8_pre_bht = _RAND_119[6:0];
  _RAND_120 = {1{`RANDOM}};
  btb_8_pre_lookup_value = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  btb_8_pre_decoder_branchD_flag = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  btb_8_pre_decoder_jump = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  btb_8_pre_decoder_branchdata = _RAND_123[5:0];
  _RAND_124 = {1{`RANDOM}};
  btb_8_pre_decoder_jr = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  btb_8_true_branch_state = _RAND_125[0:0];
  _RAND_126 = {2{`RANDOM}};
  btb_9_pc = _RAND_126[63:0];
  _RAND_127 = {1{`RANDOM}};
  btb_9_inst = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  btb_9_exception_type = _RAND_128[1:0];
  _RAND_129 = {2{`RANDOM}};
  btb_9_pre_pc_target = _RAND_129[63:0];
  _RAND_130 = {1{`RANDOM}};
  btb_9_pre_lookup_data = _RAND_130[6:0];
  _RAND_131 = {1{`RANDOM}};
  btb_9_pre_hashcode = _RAND_131[3:0];
  _RAND_132 = {1{`RANDOM}};
  btb_9_pre_pht = _RAND_132[1:0];
  _RAND_133 = {1{`RANDOM}};
  btb_9_pre_bht = _RAND_133[6:0];
  _RAND_134 = {1{`RANDOM}};
  btb_9_pre_lookup_value = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  btb_9_pre_decoder_branchD_flag = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  btb_9_pre_decoder_jump = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  btb_9_pre_decoder_branchdata = _RAND_137[5:0];
  _RAND_138 = {1{`RANDOM}};
  btb_9_pre_decoder_jr = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  btb_9_true_branch_state = _RAND_139[0:0];
  _RAND_140 = {2{`RANDOM}};
  btb_10_pc = _RAND_140[63:0];
  _RAND_141 = {1{`RANDOM}};
  btb_10_inst = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  btb_10_exception_type = _RAND_142[1:0];
  _RAND_143 = {2{`RANDOM}};
  btb_10_pre_pc_target = _RAND_143[63:0];
  _RAND_144 = {1{`RANDOM}};
  btb_10_pre_lookup_data = _RAND_144[6:0];
  _RAND_145 = {1{`RANDOM}};
  btb_10_pre_hashcode = _RAND_145[3:0];
  _RAND_146 = {1{`RANDOM}};
  btb_10_pre_pht = _RAND_146[1:0];
  _RAND_147 = {1{`RANDOM}};
  btb_10_pre_bht = _RAND_147[6:0];
  _RAND_148 = {1{`RANDOM}};
  btb_10_pre_lookup_value = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  btb_10_pre_decoder_branchD_flag = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  btb_10_pre_decoder_jump = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  btb_10_pre_decoder_branchdata = _RAND_151[5:0];
  _RAND_152 = {1{`RANDOM}};
  btb_10_pre_decoder_jr = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  btb_10_true_branch_state = _RAND_153[0:0];
  _RAND_154 = {2{`RANDOM}};
  btb_11_pc = _RAND_154[63:0];
  _RAND_155 = {1{`RANDOM}};
  btb_11_inst = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  btb_11_exception_type = _RAND_156[1:0];
  _RAND_157 = {2{`RANDOM}};
  btb_11_pre_pc_target = _RAND_157[63:0];
  _RAND_158 = {1{`RANDOM}};
  btb_11_pre_lookup_data = _RAND_158[6:0];
  _RAND_159 = {1{`RANDOM}};
  btb_11_pre_hashcode = _RAND_159[3:0];
  _RAND_160 = {1{`RANDOM}};
  btb_11_pre_pht = _RAND_160[1:0];
  _RAND_161 = {1{`RANDOM}};
  btb_11_pre_bht = _RAND_161[6:0];
  _RAND_162 = {1{`RANDOM}};
  btb_11_pre_lookup_value = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  btb_11_pre_decoder_branchD_flag = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  btb_11_pre_decoder_jump = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  btb_11_pre_decoder_branchdata = _RAND_165[5:0];
  _RAND_166 = {1{`RANDOM}};
  btb_11_pre_decoder_jr = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  btb_11_true_branch_state = _RAND_167[0:0];
  _RAND_168 = {2{`RANDOM}};
  btb_12_pc = _RAND_168[63:0];
  _RAND_169 = {1{`RANDOM}};
  btb_12_inst = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  btb_12_exception_type = _RAND_170[1:0];
  _RAND_171 = {2{`RANDOM}};
  btb_12_pre_pc_target = _RAND_171[63:0];
  _RAND_172 = {1{`RANDOM}};
  btb_12_pre_lookup_data = _RAND_172[6:0];
  _RAND_173 = {1{`RANDOM}};
  btb_12_pre_hashcode = _RAND_173[3:0];
  _RAND_174 = {1{`RANDOM}};
  btb_12_pre_pht = _RAND_174[1:0];
  _RAND_175 = {1{`RANDOM}};
  btb_12_pre_bht = _RAND_175[6:0];
  _RAND_176 = {1{`RANDOM}};
  btb_12_pre_lookup_value = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  btb_12_pre_decoder_branchD_flag = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  btb_12_pre_decoder_jump = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  btb_12_pre_decoder_branchdata = _RAND_179[5:0];
  _RAND_180 = {1{`RANDOM}};
  btb_12_pre_decoder_jr = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  btb_12_true_branch_state = _RAND_181[0:0];
  _RAND_182 = {2{`RANDOM}};
  btb_13_pc = _RAND_182[63:0];
  _RAND_183 = {1{`RANDOM}};
  btb_13_inst = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  btb_13_exception_type = _RAND_184[1:0];
  _RAND_185 = {2{`RANDOM}};
  btb_13_pre_pc_target = _RAND_185[63:0];
  _RAND_186 = {1{`RANDOM}};
  btb_13_pre_lookup_data = _RAND_186[6:0];
  _RAND_187 = {1{`RANDOM}};
  btb_13_pre_hashcode = _RAND_187[3:0];
  _RAND_188 = {1{`RANDOM}};
  btb_13_pre_pht = _RAND_188[1:0];
  _RAND_189 = {1{`RANDOM}};
  btb_13_pre_bht = _RAND_189[6:0];
  _RAND_190 = {1{`RANDOM}};
  btb_13_pre_lookup_value = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  btb_13_pre_decoder_branchD_flag = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  btb_13_pre_decoder_jump = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  btb_13_pre_decoder_branchdata = _RAND_193[5:0];
  _RAND_194 = {1{`RANDOM}};
  btb_13_pre_decoder_jr = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  btb_13_true_branch_state = _RAND_195[0:0];
  _RAND_196 = {2{`RANDOM}};
  btb_14_pc = _RAND_196[63:0];
  _RAND_197 = {1{`RANDOM}};
  btb_14_inst = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  btb_14_exception_type = _RAND_198[1:0];
  _RAND_199 = {2{`RANDOM}};
  btb_14_pre_pc_target = _RAND_199[63:0];
  _RAND_200 = {1{`RANDOM}};
  btb_14_pre_lookup_data = _RAND_200[6:0];
  _RAND_201 = {1{`RANDOM}};
  btb_14_pre_hashcode = _RAND_201[3:0];
  _RAND_202 = {1{`RANDOM}};
  btb_14_pre_pht = _RAND_202[1:0];
  _RAND_203 = {1{`RANDOM}};
  btb_14_pre_bht = _RAND_203[6:0];
  _RAND_204 = {1{`RANDOM}};
  btb_14_pre_lookup_value = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  btb_14_pre_decoder_branchD_flag = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  btb_14_pre_decoder_jump = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  btb_14_pre_decoder_branchdata = _RAND_207[5:0];
  _RAND_208 = {1{`RANDOM}};
  btb_14_pre_decoder_jr = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  btb_14_true_branch_state = _RAND_209[0:0];
  _RAND_210 = {2{`RANDOM}};
  btb_15_pc = _RAND_210[63:0];
  _RAND_211 = {1{`RANDOM}};
  btb_15_inst = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  btb_15_exception_type = _RAND_212[1:0];
  _RAND_213 = {2{`RANDOM}};
  btb_15_pre_pc_target = _RAND_213[63:0];
  _RAND_214 = {1{`RANDOM}};
  btb_15_pre_lookup_data = _RAND_214[6:0];
  _RAND_215 = {1{`RANDOM}};
  btb_15_pre_hashcode = _RAND_215[3:0];
  _RAND_216 = {1{`RANDOM}};
  btb_15_pre_pht = _RAND_216[1:0];
  _RAND_217 = {1{`RANDOM}};
  btb_15_pre_bht = _RAND_217[6:0];
  _RAND_218 = {1{`RANDOM}};
  btb_15_pre_lookup_value = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  btb_15_pre_decoder_branchD_flag = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  btb_15_pre_decoder_jump = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  btb_15_pre_decoder_branchdata = _RAND_221[5:0];
  _RAND_222 = {1{`RANDOM}};
  btb_15_pre_decoder_jr = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  btb_15_true_branch_state = _RAND_223[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    btb_0_pc = 64'h0;
  end
  if (reset) begin
    btb_0_inst = 32'h0;
  end
  if (reset) begin
    btb_0_exception_type = 2'h0;
  end
  if (reset) begin
    btb_0_pre_pc_target = 64'h0;
  end
  if (reset) begin
    btb_0_pre_lookup_data = 7'h0;
  end
  if (reset) begin
    btb_0_pre_hashcode = 4'h0;
  end
  if (reset) begin
    btb_0_pre_pht = 2'h0;
  end
  if (reset) begin
    btb_0_pre_bht = 7'h0;
  end
  if (reset) begin
    btb_0_pre_lookup_value = 8'h0;
  end
  if (reset) begin
    btb_0_pre_decoder_branchD_flag = 1'h0;
  end
  if (reset) begin
    btb_0_pre_decoder_jump = 1'h0;
  end
  if (reset) begin
    btb_0_pre_decoder_branchdata = 6'h0;
  end
  if (reset) begin
    btb_0_pre_decoder_jr = 1'h0;
  end
  if (reset) begin
    btb_0_true_branch_state = 1'h0;
  end
  if (reset) begin
    btb_1_pc = 64'h0;
  end
  if (reset) begin
    btb_1_inst = 32'h0;
  end
  if (reset) begin
    btb_1_exception_type = 2'h0;
  end
  if (reset) begin
    btb_1_pre_pc_target = 64'h0;
  end
  if (reset) begin
    btb_1_pre_lookup_data = 7'h0;
  end
  if (reset) begin
    btb_1_pre_hashcode = 4'h0;
  end
  if (reset) begin
    btb_1_pre_pht = 2'h0;
  end
  if (reset) begin
    btb_1_pre_bht = 7'h0;
  end
  if (reset) begin
    btb_1_pre_lookup_value = 8'h0;
  end
  if (reset) begin
    btb_1_pre_decoder_branchD_flag = 1'h0;
  end
  if (reset) begin
    btb_1_pre_decoder_jump = 1'h0;
  end
  if (reset) begin
    btb_1_pre_decoder_branchdata = 6'h0;
  end
  if (reset) begin
    btb_1_pre_decoder_jr = 1'h0;
  end
  if (reset) begin
    btb_1_true_branch_state = 1'h0;
  end
  if (reset) begin
    btb_2_pc = 64'h0;
  end
  if (reset) begin
    btb_2_inst = 32'h0;
  end
  if (reset) begin
    btb_2_exception_type = 2'h0;
  end
  if (reset) begin
    btb_2_pre_pc_target = 64'h0;
  end
  if (reset) begin
    btb_2_pre_lookup_data = 7'h0;
  end
  if (reset) begin
    btb_2_pre_hashcode = 4'h0;
  end
  if (reset) begin
    btb_2_pre_pht = 2'h0;
  end
  if (reset) begin
    btb_2_pre_bht = 7'h0;
  end
  if (reset) begin
    btb_2_pre_lookup_value = 8'h0;
  end
  if (reset) begin
    btb_2_pre_decoder_branchD_flag = 1'h0;
  end
  if (reset) begin
    btb_2_pre_decoder_jump = 1'h0;
  end
  if (reset) begin
    btb_2_pre_decoder_branchdata = 6'h0;
  end
  if (reset) begin
    btb_2_pre_decoder_jr = 1'h0;
  end
  if (reset) begin
    btb_2_true_branch_state = 1'h0;
  end
  if (reset) begin
    btb_3_pc = 64'h0;
  end
  if (reset) begin
    btb_3_inst = 32'h0;
  end
  if (reset) begin
    btb_3_exception_type = 2'h0;
  end
  if (reset) begin
    btb_3_pre_pc_target = 64'h0;
  end
  if (reset) begin
    btb_3_pre_lookup_data = 7'h0;
  end
  if (reset) begin
    btb_3_pre_hashcode = 4'h0;
  end
  if (reset) begin
    btb_3_pre_pht = 2'h0;
  end
  if (reset) begin
    btb_3_pre_bht = 7'h0;
  end
  if (reset) begin
    btb_3_pre_lookup_value = 8'h0;
  end
  if (reset) begin
    btb_3_pre_decoder_branchD_flag = 1'h0;
  end
  if (reset) begin
    btb_3_pre_decoder_jump = 1'h0;
  end
  if (reset) begin
    btb_3_pre_decoder_branchdata = 6'h0;
  end
  if (reset) begin
    btb_3_pre_decoder_jr = 1'h0;
  end
  if (reset) begin
    btb_3_true_branch_state = 1'h0;
  end
  if (reset) begin
    btb_4_pc = 64'h0;
  end
  if (reset) begin
    btb_4_inst = 32'h0;
  end
  if (reset) begin
    btb_4_exception_type = 2'h0;
  end
  if (reset) begin
    btb_4_pre_pc_target = 64'h0;
  end
  if (reset) begin
    btb_4_pre_lookup_data = 7'h0;
  end
  if (reset) begin
    btb_4_pre_hashcode = 4'h0;
  end
  if (reset) begin
    btb_4_pre_pht = 2'h0;
  end
  if (reset) begin
    btb_4_pre_bht = 7'h0;
  end
  if (reset) begin
    btb_4_pre_lookup_value = 8'h0;
  end
  if (reset) begin
    btb_4_pre_decoder_branchD_flag = 1'h0;
  end
  if (reset) begin
    btb_4_pre_decoder_jump = 1'h0;
  end
  if (reset) begin
    btb_4_pre_decoder_branchdata = 6'h0;
  end
  if (reset) begin
    btb_4_pre_decoder_jr = 1'h0;
  end
  if (reset) begin
    btb_4_true_branch_state = 1'h0;
  end
  if (reset) begin
    btb_5_pc = 64'h0;
  end
  if (reset) begin
    btb_5_inst = 32'h0;
  end
  if (reset) begin
    btb_5_exception_type = 2'h0;
  end
  if (reset) begin
    btb_5_pre_pc_target = 64'h0;
  end
  if (reset) begin
    btb_5_pre_lookup_data = 7'h0;
  end
  if (reset) begin
    btb_5_pre_hashcode = 4'h0;
  end
  if (reset) begin
    btb_5_pre_pht = 2'h0;
  end
  if (reset) begin
    btb_5_pre_bht = 7'h0;
  end
  if (reset) begin
    btb_5_pre_lookup_value = 8'h0;
  end
  if (reset) begin
    btb_5_pre_decoder_branchD_flag = 1'h0;
  end
  if (reset) begin
    btb_5_pre_decoder_jump = 1'h0;
  end
  if (reset) begin
    btb_5_pre_decoder_branchdata = 6'h0;
  end
  if (reset) begin
    btb_5_pre_decoder_jr = 1'h0;
  end
  if (reset) begin
    btb_5_true_branch_state = 1'h0;
  end
  if (reset) begin
    btb_6_pc = 64'h0;
  end
  if (reset) begin
    btb_6_inst = 32'h0;
  end
  if (reset) begin
    btb_6_exception_type = 2'h0;
  end
  if (reset) begin
    btb_6_pre_pc_target = 64'h0;
  end
  if (reset) begin
    btb_6_pre_lookup_data = 7'h0;
  end
  if (reset) begin
    btb_6_pre_hashcode = 4'h0;
  end
  if (reset) begin
    btb_6_pre_pht = 2'h0;
  end
  if (reset) begin
    btb_6_pre_bht = 7'h0;
  end
  if (reset) begin
    btb_6_pre_lookup_value = 8'h0;
  end
  if (reset) begin
    btb_6_pre_decoder_branchD_flag = 1'h0;
  end
  if (reset) begin
    btb_6_pre_decoder_jump = 1'h0;
  end
  if (reset) begin
    btb_6_pre_decoder_branchdata = 6'h0;
  end
  if (reset) begin
    btb_6_pre_decoder_jr = 1'h0;
  end
  if (reset) begin
    btb_6_true_branch_state = 1'h0;
  end
  if (reset) begin
    btb_7_pc = 64'h0;
  end
  if (reset) begin
    btb_7_inst = 32'h0;
  end
  if (reset) begin
    btb_7_exception_type = 2'h0;
  end
  if (reset) begin
    btb_7_pre_pc_target = 64'h0;
  end
  if (reset) begin
    btb_7_pre_lookup_data = 7'h0;
  end
  if (reset) begin
    btb_7_pre_hashcode = 4'h0;
  end
  if (reset) begin
    btb_7_pre_pht = 2'h0;
  end
  if (reset) begin
    btb_7_pre_bht = 7'h0;
  end
  if (reset) begin
    btb_7_pre_lookup_value = 8'h0;
  end
  if (reset) begin
    btb_7_pre_decoder_branchD_flag = 1'h0;
  end
  if (reset) begin
    btb_7_pre_decoder_jump = 1'h0;
  end
  if (reset) begin
    btb_7_pre_decoder_branchdata = 6'h0;
  end
  if (reset) begin
    btb_7_pre_decoder_jr = 1'h0;
  end
  if (reset) begin
    btb_7_true_branch_state = 1'h0;
  end
  if (reset) begin
    btb_8_pc = 64'h0;
  end
  if (reset) begin
    btb_8_inst = 32'h0;
  end
  if (reset) begin
    btb_8_exception_type = 2'h0;
  end
  if (reset) begin
    btb_8_pre_pc_target = 64'h0;
  end
  if (reset) begin
    btb_8_pre_lookup_data = 7'h0;
  end
  if (reset) begin
    btb_8_pre_hashcode = 4'h0;
  end
  if (reset) begin
    btb_8_pre_pht = 2'h0;
  end
  if (reset) begin
    btb_8_pre_bht = 7'h0;
  end
  if (reset) begin
    btb_8_pre_lookup_value = 8'h0;
  end
  if (reset) begin
    btb_8_pre_decoder_branchD_flag = 1'h0;
  end
  if (reset) begin
    btb_8_pre_decoder_jump = 1'h0;
  end
  if (reset) begin
    btb_8_pre_decoder_branchdata = 6'h0;
  end
  if (reset) begin
    btb_8_pre_decoder_jr = 1'h0;
  end
  if (reset) begin
    btb_8_true_branch_state = 1'h0;
  end
  if (reset) begin
    btb_9_pc = 64'h0;
  end
  if (reset) begin
    btb_9_inst = 32'h0;
  end
  if (reset) begin
    btb_9_exception_type = 2'h0;
  end
  if (reset) begin
    btb_9_pre_pc_target = 64'h0;
  end
  if (reset) begin
    btb_9_pre_lookup_data = 7'h0;
  end
  if (reset) begin
    btb_9_pre_hashcode = 4'h0;
  end
  if (reset) begin
    btb_9_pre_pht = 2'h0;
  end
  if (reset) begin
    btb_9_pre_bht = 7'h0;
  end
  if (reset) begin
    btb_9_pre_lookup_value = 8'h0;
  end
  if (reset) begin
    btb_9_pre_decoder_branchD_flag = 1'h0;
  end
  if (reset) begin
    btb_9_pre_decoder_jump = 1'h0;
  end
  if (reset) begin
    btb_9_pre_decoder_branchdata = 6'h0;
  end
  if (reset) begin
    btb_9_pre_decoder_jr = 1'h0;
  end
  if (reset) begin
    btb_9_true_branch_state = 1'h0;
  end
  if (reset) begin
    btb_10_pc = 64'h0;
  end
  if (reset) begin
    btb_10_inst = 32'h0;
  end
  if (reset) begin
    btb_10_exception_type = 2'h0;
  end
  if (reset) begin
    btb_10_pre_pc_target = 64'h0;
  end
  if (reset) begin
    btb_10_pre_lookup_data = 7'h0;
  end
  if (reset) begin
    btb_10_pre_hashcode = 4'h0;
  end
  if (reset) begin
    btb_10_pre_pht = 2'h0;
  end
  if (reset) begin
    btb_10_pre_bht = 7'h0;
  end
  if (reset) begin
    btb_10_pre_lookup_value = 8'h0;
  end
  if (reset) begin
    btb_10_pre_decoder_branchD_flag = 1'h0;
  end
  if (reset) begin
    btb_10_pre_decoder_jump = 1'h0;
  end
  if (reset) begin
    btb_10_pre_decoder_branchdata = 6'h0;
  end
  if (reset) begin
    btb_10_pre_decoder_jr = 1'h0;
  end
  if (reset) begin
    btb_10_true_branch_state = 1'h0;
  end
  if (reset) begin
    btb_11_pc = 64'h0;
  end
  if (reset) begin
    btb_11_inst = 32'h0;
  end
  if (reset) begin
    btb_11_exception_type = 2'h0;
  end
  if (reset) begin
    btb_11_pre_pc_target = 64'h0;
  end
  if (reset) begin
    btb_11_pre_lookup_data = 7'h0;
  end
  if (reset) begin
    btb_11_pre_hashcode = 4'h0;
  end
  if (reset) begin
    btb_11_pre_pht = 2'h0;
  end
  if (reset) begin
    btb_11_pre_bht = 7'h0;
  end
  if (reset) begin
    btb_11_pre_lookup_value = 8'h0;
  end
  if (reset) begin
    btb_11_pre_decoder_branchD_flag = 1'h0;
  end
  if (reset) begin
    btb_11_pre_decoder_jump = 1'h0;
  end
  if (reset) begin
    btb_11_pre_decoder_branchdata = 6'h0;
  end
  if (reset) begin
    btb_11_pre_decoder_jr = 1'h0;
  end
  if (reset) begin
    btb_11_true_branch_state = 1'h0;
  end
  if (reset) begin
    btb_12_pc = 64'h0;
  end
  if (reset) begin
    btb_12_inst = 32'h0;
  end
  if (reset) begin
    btb_12_exception_type = 2'h0;
  end
  if (reset) begin
    btb_12_pre_pc_target = 64'h0;
  end
  if (reset) begin
    btb_12_pre_lookup_data = 7'h0;
  end
  if (reset) begin
    btb_12_pre_hashcode = 4'h0;
  end
  if (reset) begin
    btb_12_pre_pht = 2'h0;
  end
  if (reset) begin
    btb_12_pre_bht = 7'h0;
  end
  if (reset) begin
    btb_12_pre_lookup_value = 8'h0;
  end
  if (reset) begin
    btb_12_pre_decoder_branchD_flag = 1'h0;
  end
  if (reset) begin
    btb_12_pre_decoder_jump = 1'h0;
  end
  if (reset) begin
    btb_12_pre_decoder_branchdata = 6'h0;
  end
  if (reset) begin
    btb_12_pre_decoder_jr = 1'h0;
  end
  if (reset) begin
    btb_12_true_branch_state = 1'h0;
  end
  if (reset) begin
    btb_13_pc = 64'h0;
  end
  if (reset) begin
    btb_13_inst = 32'h0;
  end
  if (reset) begin
    btb_13_exception_type = 2'h0;
  end
  if (reset) begin
    btb_13_pre_pc_target = 64'h0;
  end
  if (reset) begin
    btb_13_pre_lookup_data = 7'h0;
  end
  if (reset) begin
    btb_13_pre_hashcode = 4'h0;
  end
  if (reset) begin
    btb_13_pre_pht = 2'h0;
  end
  if (reset) begin
    btb_13_pre_bht = 7'h0;
  end
  if (reset) begin
    btb_13_pre_lookup_value = 8'h0;
  end
  if (reset) begin
    btb_13_pre_decoder_branchD_flag = 1'h0;
  end
  if (reset) begin
    btb_13_pre_decoder_jump = 1'h0;
  end
  if (reset) begin
    btb_13_pre_decoder_branchdata = 6'h0;
  end
  if (reset) begin
    btb_13_pre_decoder_jr = 1'h0;
  end
  if (reset) begin
    btb_13_true_branch_state = 1'h0;
  end
  if (reset) begin
    btb_14_pc = 64'h0;
  end
  if (reset) begin
    btb_14_inst = 32'h0;
  end
  if (reset) begin
    btb_14_exception_type = 2'h0;
  end
  if (reset) begin
    btb_14_pre_pc_target = 64'h0;
  end
  if (reset) begin
    btb_14_pre_lookup_data = 7'h0;
  end
  if (reset) begin
    btb_14_pre_hashcode = 4'h0;
  end
  if (reset) begin
    btb_14_pre_pht = 2'h0;
  end
  if (reset) begin
    btb_14_pre_bht = 7'h0;
  end
  if (reset) begin
    btb_14_pre_lookup_value = 8'h0;
  end
  if (reset) begin
    btb_14_pre_decoder_branchD_flag = 1'h0;
  end
  if (reset) begin
    btb_14_pre_decoder_jump = 1'h0;
  end
  if (reset) begin
    btb_14_pre_decoder_branchdata = 6'h0;
  end
  if (reset) begin
    btb_14_pre_decoder_jr = 1'h0;
  end
  if (reset) begin
    btb_14_true_branch_state = 1'h0;
  end
  if (reset) begin
    btb_15_pc = 64'h0;
  end
  if (reset) begin
    btb_15_inst = 32'h0;
  end
  if (reset) begin
    btb_15_exception_type = 2'h0;
  end
  if (reset) begin
    btb_15_pre_pc_target = 64'h0;
  end
  if (reset) begin
    btb_15_pre_lookup_data = 7'h0;
  end
  if (reset) begin
    btb_15_pre_hashcode = 4'h0;
  end
  if (reset) begin
    btb_15_pre_pht = 2'h0;
  end
  if (reset) begin
    btb_15_pre_bht = 7'h0;
  end
  if (reset) begin
    btb_15_pre_lookup_value = 8'h0;
  end
  if (reset) begin
    btb_15_pre_decoder_branchD_flag = 1'h0;
  end
  if (reset) begin
    btb_15_pre_decoder_jump = 1'h0;
  end
  if (reset) begin
    btb_15_pre_decoder_branchdata = 6'h0;
  end
  if (reset) begin
    btb_15_pre_decoder_jr = 1'h0;
  end
  if (reset) begin
    btb_15_true_branch_state = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module fifo_with_bundle(
  input         clock,
  input         reset,
  input  [1:0]  io_read_en,
  input  [1:0]  io_write_en,
  output [63:0] io_read_out_0_pc,
  output [31:0] io_read_out_0_inst,
  output [1:0]  io_read_out_0_exception_type,
  output [63:0] io_read_out_0_pre_pc_target,
  output [6:0]  io_read_out_0_pre_lookup_data,
  output [3:0]  io_read_out_0_pre_hashcode,
  output [1:0]  io_read_out_0_pre_pht,
  output [6:0]  io_read_out_0_pre_bht,
  output [7:0]  io_read_out_0_pre_lookup_value,
  output        io_read_out_0_pre_decoder_branchD_flag,
  output        io_read_out_0_pre_decoder_jump,
  output [5:0]  io_read_out_0_pre_decoder_branchdata,
  output        io_read_out_0_pre_decoder_jr,
  output        io_read_out_0_true_branch_state,
  input  [63:0] io_write_in_0_pc,
  input  [31:0] io_write_in_0_inst,
  input  [63:0] io_write_in_0_pre_pc_target,
  input  [6:0]  io_write_in_0_pre_lookup_data,
  input  [3:0]  io_write_in_0_pre_hashcode,
  input  [1:0]  io_write_in_0_pre_pht,
  input  [6:0]  io_write_in_0_pre_bht,
  input  [7:0]  io_write_in_0_pre_lookup_value,
  input         io_write_in_0_pre_decoder_branchD_flag,
  input         io_write_in_0_pre_decoder_jump,
  input  [5:0]  io_write_in_0_pre_decoder_branchdata,
  input         io_write_in_0_pre_decoder_jr,
  input         io_write_in_0_true_branch_state,
  output        io_full,
  output        io_empty,
  input         io_point_write_en,
  input         io_point_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  Look_up_table_read_first_with_bundle_clock; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_reset; // @[fifo.scala 151:55]
  wire [3:0] Look_up_table_read_first_with_bundle_io_ar_addr; // @[fifo.scala 151:55]
  wire [3:0] Look_up_table_read_first_with_bundle_io_aw_addr; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_io_write; // @[fifo.scala 151:55]
  wire [63:0] Look_up_table_read_first_with_bundle_io_in_pc; // @[fifo.scala 151:55]
  wire [31:0] Look_up_table_read_first_with_bundle_io_in_inst; // @[fifo.scala 151:55]
  wire [63:0] Look_up_table_read_first_with_bundle_io_in_pre_pc_target; // @[fifo.scala 151:55]
  wire [6:0] Look_up_table_read_first_with_bundle_io_in_pre_lookup_data; // @[fifo.scala 151:55]
  wire [3:0] Look_up_table_read_first_with_bundle_io_in_pre_hashcode; // @[fifo.scala 151:55]
  wire [1:0] Look_up_table_read_first_with_bundle_io_in_pre_pht; // @[fifo.scala 151:55]
  wire [6:0] Look_up_table_read_first_with_bundle_io_in_pre_bht; // @[fifo.scala 151:55]
  wire [7:0] Look_up_table_read_first_with_bundle_io_in_pre_lookup_value; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_io_in_pre_decoder_branchD_flag; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_io_in_pre_decoder_jump; // @[fifo.scala 151:55]
  wire [5:0] Look_up_table_read_first_with_bundle_io_in_pre_decoder_branchdata; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_io_in_pre_decoder_jr; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_io_in_true_branch_state; // @[fifo.scala 151:55]
  wire [63:0] Look_up_table_read_first_with_bundle_io_out_pc; // @[fifo.scala 151:55]
  wire [31:0] Look_up_table_read_first_with_bundle_io_out_inst; // @[fifo.scala 151:55]
  wire [1:0] Look_up_table_read_first_with_bundle_io_out_exception_type; // @[fifo.scala 151:55]
  wire [63:0] Look_up_table_read_first_with_bundle_io_out_pre_pc_target; // @[fifo.scala 151:55]
  wire [6:0] Look_up_table_read_first_with_bundle_io_out_pre_lookup_data; // @[fifo.scala 151:55]
  wire [3:0] Look_up_table_read_first_with_bundle_io_out_pre_hashcode; // @[fifo.scala 151:55]
  wire [1:0] Look_up_table_read_first_with_bundle_io_out_pre_pht; // @[fifo.scala 151:55]
  wire [6:0] Look_up_table_read_first_with_bundle_io_out_pre_bht; // @[fifo.scala 151:55]
  wire [7:0] Look_up_table_read_first_with_bundle_io_out_pre_lookup_value; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_io_out_pre_decoder_branchD_flag; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_io_out_pre_decoder_jump; // @[fifo.scala 151:55]
  wire [5:0] Look_up_table_read_first_with_bundle_io_out_pre_decoder_branchdata; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_io_out_pre_decoder_jr; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_io_out_true_branch_state; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_1_clock; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_1_reset; // @[fifo.scala 151:55]
  wire [3:0] Look_up_table_read_first_with_bundle_1_io_ar_addr; // @[fifo.scala 151:55]
  wire [3:0] Look_up_table_read_first_with_bundle_1_io_aw_addr; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_1_io_write; // @[fifo.scala 151:55]
  wire [63:0] Look_up_table_read_first_with_bundle_1_io_in_pc; // @[fifo.scala 151:55]
  wire [31:0] Look_up_table_read_first_with_bundle_1_io_in_inst; // @[fifo.scala 151:55]
  wire [63:0] Look_up_table_read_first_with_bundle_1_io_in_pre_pc_target; // @[fifo.scala 151:55]
  wire [6:0] Look_up_table_read_first_with_bundle_1_io_in_pre_lookup_data; // @[fifo.scala 151:55]
  wire [3:0] Look_up_table_read_first_with_bundle_1_io_in_pre_hashcode; // @[fifo.scala 151:55]
  wire [1:0] Look_up_table_read_first_with_bundle_1_io_in_pre_pht; // @[fifo.scala 151:55]
  wire [6:0] Look_up_table_read_first_with_bundle_1_io_in_pre_bht; // @[fifo.scala 151:55]
  wire [7:0] Look_up_table_read_first_with_bundle_1_io_in_pre_lookup_value; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_1_io_in_pre_decoder_branchD_flag; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_1_io_in_pre_decoder_jump; // @[fifo.scala 151:55]
  wire [5:0] Look_up_table_read_first_with_bundle_1_io_in_pre_decoder_branchdata; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_1_io_in_pre_decoder_jr; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_1_io_in_true_branch_state; // @[fifo.scala 151:55]
  wire [63:0] Look_up_table_read_first_with_bundle_1_io_out_pc; // @[fifo.scala 151:55]
  wire [31:0] Look_up_table_read_first_with_bundle_1_io_out_inst; // @[fifo.scala 151:55]
  wire [1:0] Look_up_table_read_first_with_bundle_1_io_out_exception_type; // @[fifo.scala 151:55]
  wire [63:0] Look_up_table_read_first_with_bundle_1_io_out_pre_pc_target; // @[fifo.scala 151:55]
  wire [6:0] Look_up_table_read_first_with_bundle_1_io_out_pre_lookup_data; // @[fifo.scala 151:55]
  wire [3:0] Look_up_table_read_first_with_bundle_1_io_out_pre_hashcode; // @[fifo.scala 151:55]
  wire [1:0] Look_up_table_read_first_with_bundle_1_io_out_pre_pht; // @[fifo.scala 151:55]
  wire [6:0] Look_up_table_read_first_with_bundle_1_io_out_pre_bht; // @[fifo.scala 151:55]
  wire [7:0] Look_up_table_read_first_with_bundle_1_io_out_pre_lookup_value; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_1_io_out_pre_decoder_branchD_flag; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_1_io_out_pre_decoder_jump; // @[fifo.scala 151:55]
  wire [5:0] Look_up_table_read_first_with_bundle_1_io_out_pre_decoder_branchdata; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_1_io_out_pre_decoder_jr; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_1_io_out_true_branch_state; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_2_clock; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_2_reset; // @[fifo.scala 151:55]
  wire [3:0] Look_up_table_read_first_with_bundle_2_io_ar_addr; // @[fifo.scala 151:55]
  wire [3:0] Look_up_table_read_first_with_bundle_2_io_aw_addr; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_2_io_write; // @[fifo.scala 151:55]
  wire [63:0] Look_up_table_read_first_with_bundle_2_io_in_pc; // @[fifo.scala 151:55]
  wire [31:0] Look_up_table_read_first_with_bundle_2_io_in_inst; // @[fifo.scala 151:55]
  wire [63:0] Look_up_table_read_first_with_bundle_2_io_in_pre_pc_target; // @[fifo.scala 151:55]
  wire [6:0] Look_up_table_read_first_with_bundle_2_io_in_pre_lookup_data; // @[fifo.scala 151:55]
  wire [3:0] Look_up_table_read_first_with_bundle_2_io_in_pre_hashcode; // @[fifo.scala 151:55]
  wire [1:0] Look_up_table_read_first_with_bundle_2_io_in_pre_pht; // @[fifo.scala 151:55]
  wire [6:0] Look_up_table_read_first_with_bundle_2_io_in_pre_bht; // @[fifo.scala 151:55]
  wire [7:0] Look_up_table_read_first_with_bundle_2_io_in_pre_lookup_value; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_2_io_in_pre_decoder_branchD_flag; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_2_io_in_pre_decoder_jump; // @[fifo.scala 151:55]
  wire [5:0] Look_up_table_read_first_with_bundle_2_io_in_pre_decoder_branchdata; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_2_io_in_pre_decoder_jr; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_2_io_in_true_branch_state; // @[fifo.scala 151:55]
  wire [63:0] Look_up_table_read_first_with_bundle_2_io_out_pc; // @[fifo.scala 151:55]
  wire [31:0] Look_up_table_read_first_with_bundle_2_io_out_inst; // @[fifo.scala 151:55]
  wire [1:0] Look_up_table_read_first_with_bundle_2_io_out_exception_type; // @[fifo.scala 151:55]
  wire [63:0] Look_up_table_read_first_with_bundle_2_io_out_pre_pc_target; // @[fifo.scala 151:55]
  wire [6:0] Look_up_table_read_first_with_bundle_2_io_out_pre_lookup_data; // @[fifo.scala 151:55]
  wire [3:0] Look_up_table_read_first_with_bundle_2_io_out_pre_hashcode; // @[fifo.scala 151:55]
  wire [1:0] Look_up_table_read_first_with_bundle_2_io_out_pre_pht; // @[fifo.scala 151:55]
  wire [6:0] Look_up_table_read_first_with_bundle_2_io_out_pre_bht; // @[fifo.scala 151:55]
  wire [7:0] Look_up_table_read_first_with_bundle_2_io_out_pre_lookup_value; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_2_io_out_pre_decoder_branchD_flag; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_2_io_out_pre_decoder_jump; // @[fifo.scala 151:55]
  wire [5:0] Look_up_table_read_first_with_bundle_2_io_out_pre_decoder_branchdata; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_2_io_out_pre_decoder_jr; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_2_io_out_true_branch_state; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_3_clock; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_3_reset; // @[fifo.scala 151:55]
  wire [3:0] Look_up_table_read_first_with_bundle_3_io_ar_addr; // @[fifo.scala 151:55]
  wire [3:0] Look_up_table_read_first_with_bundle_3_io_aw_addr; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_3_io_write; // @[fifo.scala 151:55]
  wire [63:0] Look_up_table_read_first_with_bundle_3_io_in_pc; // @[fifo.scala 151:55]
  wire [31:0] Look_up_table_read_first_with_bundle_3_io_in_inst; // @[fifo.scala 151:55]
  wire [63:0] Look_up_table_read_first_with_bundle_3_io_in_pre_pc_target; // @[fifo.scala 151:55]
  wire [6:0] Look_up_table_read_first_with_bundle_3_io_in_pre_lookup_data; // @[fifo.scala 151:55]
  wire [3:0] Look_up_table_read_first_with_bundle_3_io_in_pre_hashcode; // @[fifo.scala 151:55]
  wire [1:0] Look_up_table_read_first_with_bundle_3_io_in_pre_pht; // @[fifo.scala 151:55]
  wire [6:0] Look_up_table_read_first_with_bundle_3_io_in_pre_bht; // @[fifo.scala 151:55]
  wire [7:0] Look_up_table_read_first_with_bundle_3_io_in_pre_lookup_value; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_3_io_in_pre_decoder_branchD_flag; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_3_io_in_pre_decoder_jump; // @[fifo.scala 151:55]
  wire [5:0] Look_up_table_read_first_with_bundle_3_io_in_pre_decoder_branchdata; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_3_io_in_pre_decoder_jr; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_3_io_in_true_branch_state; // @[fifo.scala 151:55]
  wire [63:0] Look_up_table_read_first_with_bundle_3_io_out_pc; // @[fifo.scala 151:55]
  wire [31:0] Look_up_table_read_first_with_bundle_3_io_out_inst; // @[fifo.scala 151:55]
  wire [1:0] Look_up_table_read_first_with_bundle_3_io_out_exception_type; // @[fifo.scala 151:55]
  wire [63:0] Look_up_table_read_first_with_bundle_3_io_out_pre_pc_target; // @[fifo.scala 151:55]
  wire [6:0] Look_up_table_read_first_with_bundle_3_io_out_pre_lookup_data; // @[fifo.scala 151:55]
  wire [3:0] Look_up_table_read_first_with_bundle_3_io_out_pre_hashcode; // @[fifo.scala 151:55]
  wire [1:0] Look_up_table_read_first_with_bundle_3_io_out_pre_pht; // @[fifo.scala 151:55]
  wire [6:0] Look_up_table_read_first_with_bundle_3_io_out_pre_bht; // @[fifo.scala 151:55]
  wire [7:0] Look_up_table_read_first_with_bundle_3_io_out_pre_lookup_value; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_3_io_out_pre_decoder_branchD_flag; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_3_io_out_pre_decoder_jump; // @[fifo.scala 151:55]
  wire [5:0] Look_up_table_read_first_with_bundle_3_io_out_pre_decoder_branchdata; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_3_io_out_pre_decoder_jr; // @[fifo.scala 151:55]
  wire  Look_up_table_read_first_with_bundle_3_io_out_true_branch_state; // @[fifo.scala 151:55]
  reg [1:0] write_banks_points; // @[fifo.scala 152:37]
  reg [3:0] write_length_points; // @[fifo.scala 153:38]
  reg [1:0] read_banks_points; // @[fifo.scala 154:36]
  reg [3:0] read_length_points; // @[fifo.scala 155:37]
  wire  _fifo_banks_3_write_T_1 = write_banks_points == 2'h3; // @[Mux.scala 81:61]
  wire  _write_banks_points_T = io_point_flush | io_point_write_en; // @[fifo.scala 175:46]
  wire [1:0] _write_banks_points_T_2 = write_banks_points + io_write_en; // @[fifo.scala 175:91]
  wire [2:0] _write_length_points_T_1 = {1'h0,write_banks_points}; // @[Cat.scala 31:58]
  wire [2:0] _GEN_56 = {{1'd0}, io_write_en}; // @[fifo.scala 176:134]
  wire [2:0] _write_length_points_T_3 = _write_length_points_T_1 + _GEN_56; // @[fifo.scala 176:134]
  wire [3:0] _GEN_57 = {{3'd0}, _write_length_points_T_3[2]}; // @[fifo.scala 176:93]
  wire [3:0] _write_length_points_T_7 = write_length_points + _GEN_57; // @[fifo.scala 176:93]
  wire [1:0] _read_banks_points_T_2 = read_banks_points + io_read_en; // @[fifo.scala 177:89]
  wire [2:0] _read_length_points_T_1 = {1'h0,read_banks_points}; // @[Cat.scala 31:58]
  wire [2:0] _GEN_58 = {{1'd0}, io_read_en}; // @[fifo.scala 178:131]
  wire [2:0] _read_length_points_T_3 = _read_length_points_T_1 + _GEN_58; // @[fifo.scala 178:131]
  wire [3:0] _GEN_59 = {{3'd0}, _read_length_points_T_3[2]}; // @[fifo.scala 178:92]
  wire [3:0] _read_length_points_T_7 = read_length_points + _GEN_59; // @[fifo.scala 178:92]
  wire [63:0] fifo_banks_0_out_pc = Look_up_table_read_first_with_bundle_io_out_pc; // @[fifo.scala 151:{29,29}]
  wire [31:0] fifo_banks_0_out_inst = Look_up_table_read_first_with_bundle_io_out_inst; // @[fifo.scala 151:{29,29}]
  wire [1:0] fifo_banks_0_out_exception_type = Look_up_table_read_first_with_bundle_io_out_exception_type; // @[fifo.scala 151:{29,29}]
  wire [63:0] fifo_banks_0_out_pre_pc_target = Look_up_table_read_first_with_bundle_io_out_pre_pc_target; // @[fifo.scala 151:{29,29}]
  wire [6:0] fifo_banks_0_out_pre_lookup_data = Look_up_table_read_first_with_bundle_io_out_pre_lookup_data; // @[fifo.scala 151:{29,29}]
  wire [3:0] fifo_banks_0_out_pre_hashcode = Look_up_table_read_first_with_bundle_io_out_pre_hashcode; // @[fifo.scala 151:{29,29}]
  wire [1:0] fifo_banks_0_out_pre_pht = Look_up_table_read_first_with_bundle_io_out_pre_pht; // @[fifo.scala 151:{29,29}]
  wire [6:0] fifo_banks_0_out_pre_bht = Look_up_table_read_first_with_bundle_io_out_pre_bht; // @[fifo.scala 151:{29,29}]
  wire [7:0] fifo_banks_0_out_pre_lookup_value = Look_up_table_read_first_with_bundle_io_out_pre_lookup_value; // @[fifo.scala 151:{29,29}]
  wire  fifo_banks_0_out_pre_decoder_branchD_flag = Look_up_table_read_first_with_bundle_io_out_pre_decoder_branchD_flag
    ; // @[fifo.scala 151:{29,29}]
  wire  fifo_banks_0_out_pre_decoder_jump = Look_up_table_read_first_with_bundle_io_out_pre_decoder_jump; // @[fifo.scala 151:{29,29}]
  wire [5:0] fifo_banks_0_out_pre_decoder_branchdata =
    Look_up_table_read_first_with_bundle_io_out_pre_decoder_branchdata; // @[fifo.scala 151:{29,29}]
  wire  fifo_banks_0_out_pre_decoder_jr = Look_up_table_read_first_with_bundle_io_out_pre_decoder_jr; // @[fifo.scala 151:{29,29}]
  wire  fifo_banks_0_out_true_branch_state = Look_up_table_read_first_with_bundle_io_out_true_branch_state; // @[fifo.scala 151:{29,29}]
  wire [63:0] fifo_banks_1_out_pc = Look_up_table_read_first_with_bundle_1_io_out_pc; // @[fifo.scala 151:{29,29}]
  wire [63:0] _GEN_14 = 2'h1 == read_banks_points ? fifo_banks_1_out_pc : fifo_banks_0_out_pc; // @[fifo.scala 180:{30,30}]
  wire [31:0] fifo_banks_1_out_inst = Look_up_table_read_first_with_bundle_1_io_out_inst; // @[fifo.scala 151:{29,29}]
  wire [31:0] _GEN_15 = 2'h1 == read_banks_points ? fifo_banks_1_out_inst : fifo_banks_0_out_inst; // @[fifo.scala 180:{30,30}]
  wire [1:0] fifo_banks_1_out_exception_type = Look_up_table_read_first_with_bundle_1_io_out_exception_type; // @[fifo.scala 151:{29,29}]
  wire [1:0] _GEN_16 = 2'h1 == read_banks_points ? fifo_banks_1_out_exception_type : fifo_banks_0_out_exception_type; // @[fifo.scala 180:{30,30}]
  wire [63:0] fifo_banks_1_out_pre_pc_target = Look_up_table_read_first_with_bundle_1_io_out_pre_pc_target; // @[fifo.scala 151:{29,29}]
  wire [63:0] _GEN_17 = 2'h1 == read_banks_points ? fifo_banks_1_out_pre_pc_target : fifo_banks_0_out_pre_pc_target; // @[fifo.scala 180:{30,30}]
  wire [6:0] fifo_banks_1_out_pre_lookup_data = Look_up_table_read_first_with_bundle_1_io_out_pre_lookup_data; // @[fifo.scala 151:{29,29}]
  wire [6:0] _GEN_18 = 2'h1 == read_banks_points ? fifo_banks_1_out_pre_lookup_data : fifo_banks_0_out_pre_lookup_data; // @[fifo.scala 180:{30,30}]
  wire [3:0] fifo_banks_1_out_pre_hashcode = Look_up_table_read_first_with_bundle_1_io_out_pre_hashcode; // @[fifo.scala 151:{29,29}]
  wire [3:0] _GEN_19 = 2'h1 == read_banks_points ? fifo_banks_1_out_pre_hashcode : fifo_banks_0_out_pre_hashcode; // @[fifo.scala 180:{30,30}]
  wire [1:0] fifo_banks_1_out_pre_pht = Look_up_table_read_first_with_bundle_1_io_out_pre_pht; // @[fifo.scala 151:{29,29}]
  wire [1:0] _GEN_20 = 2'h1 == read_banks_points ? fifo_banks_1_out_pre_pht : fifo_banks_0_out_pre_pht; // @[fifo.scala 180:{30,30}]
  wire [6:0] fifo_banks_1_out_pre_bht = Look_up_table_read_first_with_bundle_1_io_out_pre_bht; // @[fifo.scala 151:{29,29}]
  wire [6:0] _GEN_21 = 2'h1 == read_banks_points ? fifo_banks_1_out_pre_bht : fifo_banks_0_out_pre_bht; // @[fifo.scala 180:{30,30}]
  wire [7:0] fifo_banks_1_out_pre_lookup_value = Look_up_table_read_first_with_bundle_1_io_out_pre_lookup_value; // @[fifo.scala 151:{29,29}]
  wire [7:0] _GEN_22 = 2'h1 == read_banks_points ? fifo_banks_1_out_pre_lookup_value : fifo_banks_0_out_pre_lookup_value
    ; // @[fifo.scala 180:{30,30}]
  wire  fifo_banks_1_out_pre_decoder_branchD_flag =
    Look_up_table_read_first_with_bundle_1_io_out_pre_decoder_branchD_flag; // @[fifo.scala 151:{29,29}]
  wire  _GEN_23 = 2'h1 == read_banks_points ? fifo_banks_1_out_pre_decoder_branchD_flag :
    fifo_banks_0_out_pre_decoder_branchD_flag; // @[fifo.scala 180:{30,30}]
  wire  fifo_banks_1_out_pre_decoder_jump = Look_up_table_read_first_with_bundle_1_io_out_pre_decoder_jump; // @[fifo.scala 151:{29,29}]
  wire  _GEN_24 = 2'h1 == read_banks_points ? fifo_banks_1_out_pre_decoder_jump : fifo_banks_0_out_pre_decoder_jump; // @[fifo.scala 180:{30,30}]
  wire [5:0] fifo_banks_1_out_pre_decoder_branchdata =
    Look_up_table_read_first_with_bundle_1_io_out_pre_decoder_branchdata; // @[fifo.scala 151:{29,29}]
  wire [5:0] _GEN_25 = 2'h1 == read_banks_points ? fifo_banks_1_out_pre_decoder_branchdata :
    fifo_banks_0_out_pre_decoder_branchdata; // @[fifo.scala 180:{30,30}]
  wire  fifo_banks_1_out_pre_decoder_jr = Look_up_table_read_first_with_bundle_1_io_out_pre_decoder_jr; // @[fifo.scala 151:{29,29}]
  wire  _GEN_26 = 2'h1 == read_banks_points ? fifo_banks_1_out_pre_decoder_jr : fifo_banks_0_out_pre_decoder_jr; // @[fifo.scala 180:{30,30}]
  wire  fifo_banks_1_out_true_branch_state = Look_up_table_read_first_with_bundle_1_io_out_true_branch_state; // @[fifo.scala 151:{29,29}]
  wire  _GEN_27 = 2'h1 == read_banks_points ? fifo_banks_1_out_true_branch_state : fifo_banks_0_out_true_branch_state; // @[fifo.scala 180:{30,30}]
  wire [63:0] fifo_banks_2_out_pc = Look_up_table_read_first_with_bundle_2_io_out_pc; // @[fifo.scala 151:{29,29}]
  wire [63:0] _GEN_28 = 2'h2 == read_banks_points ? fifo_banks_2_out_pc : _GEN_14; // @[fifo.scala 180:{30,30}]
  wire [31:0] fifo_banks_2_out_inst = Look_up_table_read_first_with_bundle_2_io_out_inst; // @[fifo.scala 151:{29,29}]
  wire [31:0] _GEN_29 = 2'h2 == read_banks_points ? fifo_banks_2_out_inst : _GEN_15; // @[fifo.scala 180:{30,30}]
  wire [1:0] fifo_banks_2_out_exception_type = Look_up_table_read_first_with_bundle_2_io_out_exception_type; // @[fifo.scala 151:{29,29}]
  wire [1:0] _GEN_30 = 2'h2 == read_banks_points ? fifo_banks_2_out_exception_type : _GEN_16; // @[fifo.scala 180:{30,30}]
  wire [63:0] fifo_banks_2_out_pre_pc_target = Look_up_table_read_first_with_bundle_2_io_out_pre_pc_target; // @[fifo.scala 151:{29,29}]
  wire [63:0] _GEN_31 = 2'h2 == read_banks_points ? fifo_banks_2_out_pre_pc_target : _GEN_17; // @[fifo.scala 180:{30,30}]
  wire [6:0] fifo_banks_2_out_pre_lookup_data = Look_up_table_read_first_with_bundle_2_io_out_pre_lookup_data; // @[fifo.scala 151:{29,29}]
  wire [6:0] _GEN_32 = 2'h2 == read_banks_points ? fifo_banks_2_out_pre_lookup_data : _GEN_18; // @[fifo.scala 180:{30,30}]
  wire [3:0] fifo_banks_2_out_pre_hashcode = Look_up_table_read_first_with_bundle_2_io_out_pre_hashcode; // @[fifo.scala 151:{29,29}]
  wire [3:0] _GEN_33 = 2'h2 == read_banks_points ? fifo_banks_2_out_pre_hashcode : _GEN_19; // @[fifo.scala 180:{30,30}]
  wire [1:0] fifo_banks_2_out_pre_pht = Look_up_table_read_first_with_bundle_2_io_out_pre_pht; // @[fifo.scala 151:{29,29}]
  wire [1:0] _GEN_34 = 2'h2 == read_banks_points ? fifo_banks_2_out_pre_pht : _GEN_20; // @[fifo.scala 180:{30,30}]
  wire [6:0] fifo_banks_2_out_pre_bht = Look_up_table_read_first_with_bundle_2_io_out_pre_bht; // @[fifo.scala 151:{29,29}]
  wire [6:0] _GEN_35 = 2'h2 == read_banks_points ? fifo_banks_2_out_pre_bht : _GEN_21; // @[fifo.scala 180:{30,30}]
  wire [7:0] fifo_banks_2_out_pre_lookup_value = Look_up_table_read_first_with_bundle_2_io_out_pre_lookup_value; // @[fifo.scala 151:{29,29}]
  wire [7:0] _GEN_36 = 2'h2 == read_banks_points ? fifo_banks_2_out_pre_lookup_value : _GEN_22; // @[fifo.scala 180:{30,30}]
  wire  fifo_banks_2_out_pre_decoder_branchD_flag =
    Look_up_table_read_first_with_bundle_2_io_out_pre_decoder_branchD_flag; // @[fifo.scala 151:{29,29}]
  wire  _GEN_37 = 2'h2 == read_banks_points ? fifo_banks_2_out_pre_decoder_branchD_flag : _GEN_23; // @[fifo.scala 180:{30,30}]
  wire  fifo_banks_2_out_pre_decoder_jump = Look_up_table_read_first_with_bundle_2_io_out_pre_decoder_jump; // @[fifo.scala 151:{29,29}]
  wire  _GEN_38 = 2'h2 == read_banks_points ? fifo_banks_2_out_pre_decoder_jump : _GEN_24; // @[fifo.scala 180:{30,30}]
  wire [5:0] fifo_banks_2_out_pre_decoder_branchdata =
    Look_up_table_read_first_with_bundle_2_io_out_pre_decoder_branchdata; // @[fifo.scala 151:{29,29}]
  wire [5:0] _GEN_39 = 2'h2 == read_banks_points ? fifo_banks_2_out_pre_decoder_branchdata : _GEN_25; // @[fifo.scala 180:{30,30}]
  wire  fifo_banks_2_out_pre_decoder_jr = Look_up_table_read_first_with_bundle_2_io_out_pre_decoder_jr; // @[fifo.scala 151:{29,29}]
  wire  _GEN_40 = 2'h2 == read_banks_points ? fifo_banks_2_out_pre_decoder_jr : _GEN_26; // @[fifo.scala 180:{30,30}]
  wire  fifo_banks_2_out_true_branch_state = Look_up_table_read_first_with_bundle_2_io_out_true_branch_state; // @[fifo.scala 151:{29,29}]
  wire  _GEN_41 = 2'h2 == read_banks_points ? fifo_banks_2_out_true_branch_state : _GEN_27; // @[fifo.scala 180:{30,30}]
  wire [63:0] fifo_banks_3_out_pc = Look_up_table_read_first_with_bundle_3_io_out_pc; // @[fifo.scala 151:{29,29}]
  wire [63:0] _GEN_42 = 2'h3 == read_banks_points ? fifo_banks_3_out_pc : _GEN_28; // @[fifo.scala 180:{30,30}]
  wire [31:0] fifo_banks_3_out_inst = Look_up_table_read_first_with_bundle_3_io_out_inst; // @[fifo.scala 151:{29,29}]
  wire [31:0] _GEN_43 = 2'h3 == read_banks_points ? fifo_banks_3_out_inst : _GEN_29; // @[fifo.scala 180:{30,30}]
  wire [1:0] fifo_banks_3_out_exception_type = Look_up_table_read_first_with_bundle_3_io_out_exception_type; // @[fifo.scala 151:{29,29}]
  wire [1:0] _GEN_44 = 2'h3 == read_banks_points ? fifo_banks_3_out_exception_type : _GEN_30; // @[fifo.scala 180:{30,30}]
  wire [63:0] fifo_banks_3_out_pre_pc_target = Look_up_table_read_first_with_bundle_3_io_out_pre_pc_target; // @[fifo.scala 151:{29,29}]
  wire [63:0] _GEN_45 = 2'h3 == read_banks_points ? fifo_banks_3_out_pre_pc_target : _GEN_31; // @[fifo.scala 180:{30,30}]
  wire [6:0] fifo_banks_3_out_pre_lookup_data = Look_up_table_read_first_with_bundle_3_io_out_pre_lookup_data; // @[fifo.scala 151:{29,29}]
  wire [6:0] _GEN_46 = 2'h3 == read_banks_points ? fifo_banks_3_out_pre_lookup_data : _GEN_32; // @[fifo.scala 180:{30,30}]
  wire [3:0] fifo_banks_3_out_pre_hashcode = Look_up_table_read_first_with_bundle_3_io_out_pre_hashcode; // @[fifo.scala 151:{29,29}]
  wire [3:0] _GEN_47 = 2'h3 == read_banks_points ? fifo_banks_3_out_pre_hashcode : _GEN_33; // @[fifo.scala 180:{30,30}]
  wire [1:0] fifo_banks_3_out_pre_pht = Look_up_table_read_first_with_bundle_3_io_out_pre_pht; // @[fifo.scala 151:{29,29}]
  wire [1:0] _GEN_48 = 2'h3 == read_banks_points ? fifo_banks_3_out_pre_pht : _GEN_34; // @[fifo.scala 180:{30,30}]
  wire [6:0] fifo_banks_3_out_pre_bht = Look_up_table_read_first_with_bundle_3_io_out_pre_bht; // @[fifo.scala 151:{29,29}]
  wire [6:0] _GEN_49 = 2'h3 == read_banks_points ? fifo_banks_3_out_pre_bht : _GEN_35; // @[fifo.scala 180:{30,30}]
  wire [7:0] fifo_banks_3_out_pre_lookup_value = Look_up_table_read_first_with_bundle_3_io_out_pre_lookup_value; // @[fifo.scala 151:{29,29}]
  wire [7:0] _GEN_50 = 2'h3 == read_banks_points ? fifo_banks_3_out_pre_lookup_value : _GEN_36; // @[fifo.scala 180:{30,30}]
  wire  fifo_banks_3_out_pre_decoder_branchD_flag =
    Look_up_table_read_first_with_bundle_3_io_out_pre_decoder_branchD_flag; // @[fifo.scala 151:{29,29}]
  wire  _GEN_51 = 2'h3 == read_banks_points ? fifo_banks_3_out_pre_decoder_branchD_flag : _GEN_37; // @[fifo.scala 180:{30,30}]
  wire  fifo_banks_3_out_pre_decoder_jump = Look_up_table_read_first_with_bundle_3_io_out_pre_decoder_jump; // @[fifo.scala 151:{29,29}]
  wire  _GEN_52 = 2'h3 == read_banks_points ? fifo_banks_3_out_pre_decoder_jump : _GEN_38; // @[fifo.scala 180:{30,30}]
  wire [5:0] fifo_banks_3_out_pre_decoder_branchdata =
    Look_up_table_read_first_with_bundle_3_io_out_pre_decoder_branchdata; // @[fifo.scala 151:{29,29}]
  wire [5:0] _GEN_53 = 2'h3 == read_banks_points ? fifo_banks_3_out_pre_decoder_branchdata : _GEN_39; // @[fifo.scala 180:{30,30}]
  wire  fifo_banks_3_out_pre_decoder_jr = Look_up_table_read_first_with_bundle_3_io_out_pre_decoder_jr; // @[fifo.scala 151:{29,29}]
  wire  _GEN_54 = 2'h3 == read_banks_points ? fifo_banks_3_out_pre_decoder_jr : _GEN_40; // @[fifo.scala 180:{30,30}]
  wire  fifo_banks_3_out_true_branch_state = Look_up_table_read_first_with_bundle_3_io_out_true_branch_state; // @[fifo.scala 151:{29,29}]
  wire  _GEN_55 = 2'h3 == read_banks_points ? fifo_banks_3_out_true_branch_state : _GEN_41; // @[fifo.scala 180:{30,30}]
  wire  _io_empty_T_1 = write_length_points == read_length_points; // @[fifo.scala 187:82]
  wire [2:0] _io_full_T_3 = _write_length_points_T_1 + 3'h1; // @[fifo.scala 189:98]
  wire [3:0] _io_full_T_7 = write_length_points + 4'h1; // @[fifo.scala 190:33]
  wire  _io_full_T_12 = _io_full_T_7 == read_length_points & (_fifo_banks_3_write_T_1 & read_banks_points == 2'h0); // @[fifo.scala 190:12]
  Look_up_table_read_first_with_bundle Look_up_table_read_first_with_bundle ( // @[fifo.scala 151:55]
    .clock(Look_up_table_read_first_with_bundle_clock),
    .reset(Look_up_table_read_first_with_bundle_reset),
    .io_ar_addr(Look_up_table_read_first_with_bundle_io_ar_addr),
    .io_aw_addr(Look_up_table_read_first_with_bundle_io_aw_addr),
    .io_write(Look_up_table_read_first_with_bundle_io_write),
    .io_in_pc(Look_up_table_read_first_with_bundle_io_in_pc),
    .io_in_inst(Look_up_table_read_first_with_bundle_io_in_inst),
    .io_in_pre_pc_target(Look_up_table_read_first_with_bundle_io_in_pre_pc_target),
    .io_in_pre_lookup_data(Look_up_table_read_first_with_bundle_io_in_pre_lookup_data),
    .io_in_pre_hashcode(Look_up_table_read_first_with_bundle_io_in_pre_hashcode),
    .io_in_pre_pht(Look_up_table_read_first_with_bundle_io_in_pre_pht),
    .io_in_pre_bht(Look_up_table_read_first_with_bundle_io_in_pre_bht),
    .io_in_pre_lookup_value(Look_up_table_read_first_with_bundle_io_in_pre_lookup_value),
    .io_in_pre_decoder_branchD_flag(Look_up_table_read_first_with_bundle_io_in_pre_decoder_branchD_flag),
    .io_in_pre_decoder_jump(Look_up_table_read_first_with_bundle_io_in_pre_decoder_jump),
    .io_in_pre_decoder_branchdata(Look_up_table_read_first_with_bundle_io_in_pre_decoder_branchdata),
    .io_in_pre_decoder_jr(Look_up_table_read_first_with_bundle_io_in_pre_decoder_jr),
    .io_in_true_branch_state(Look_up_table_read_first_with_bundle_io_in_true_branch_state),
    .io_out_pc(Look_up_table_read_first_with_bundle_io_out_pc),
    .io_out_inst(Look_up_table_read_first_with_bundle_io_out_inst),
    .io_out_exception_type(Look_up_table_read_first_with_bundle_io_out_exception_type),
    .io_out_pre_pc_target(Look_up_table_read_first_with_bundle_io_out_pre_pc_target),
    .io_out_pre_lookup_data(Look_up_table_read_first_with_bundle_io_out_pre_lookup_data),
    .io_out_pre_hashcode(Look_up_table_read_first_with_bundle_io_out_pre_hashcode),
    .io_out_pre_pht(Look_up_table_read_first_with_bundle_io_out_pre_pht),
    .io_out_pre_bht(Look_up_table_read_first_with_bundle_io_out_pre_bht),
    .io_out_pre_lookup_value(Look_up_table_read_first_with_bundle_io_out_pre_lookup_value),
    .io_out_pre_decoder_branchD_flag(Look_up_table_read_first_with_bundle_io_out_pre_decoder_branchD_flag),
    .io_out_pre_decoder_jump(Look_up_table_read_first_with_bundle_io_out_pre_decoder_jump),
    .io_out_pre_decoder_branchdata(Look_up_table_read_first_with_bundle_io_out_pre_decoder_branchdata),
    .io_out_pre_decoder_jr(Look_up_table_read_first_with_bundle_io_out_pre_decoder_jr),
    .io_out_true_branch_state(Look_up_table_read_first_with_bundle_io_out_true_branch_state)
  );
  Look_up_table_read_first_with_bundle Look_up_table_read_first_with_bundle_1 ( // @[fifo.scala 151:55]
    .clock(Look_up_table_read_first_with_bundle_1_clock),
    .reset(Look_up_table_read_first_with_bundle_1_reset),
    .io_ar_addr(Look_up_table_read_first_with_bundle_1_io_ar_addr),
    .io_aw_addr(Look_up_table_read_first_with_bundle_1_io_aw_addr),
    .io_write(Look_up_table_read_first_with_bundle_1_io_write),
    .io_in_pc(Look_up_table_read_first_with_bundle_1_io_in_pc),
    .io_in_inst(Look_up_table_read_first_with_bundle_1_io_in_inst),
    .io_in_pre_pc_target(Look_up_table_read_first_with_bundle_1_io_in_pre_pc_target),
    .io_in_pre_lookup_data(Look_up_table_read_first_with_bundle_1_io_in_pre_lookup_data),
    .io_in_pre_hashcode(Look_up_table_read_first_with_bundle_1_io_in_pre_hashcode),
    .io_in_pre_pht(Look_up_table_read_first_with_bundle_1_io_in_pre_pht),
    .io_in_pre_bht(Look_up_table_read_first_with_bundle_1_io_in_pre_bht),
    .io_in_pre_lookup_value(Look_up_table_read_first_with_bundle_1_io_in_pre_lookup_value),
    .io_in_pre_decoder_branchD_flag(Look_up_table_read_first_with_bundle_1_io_in_pre_decoder_branchD_flag),
    .io_in_pre_decoder_jump(Look_up_table_read_first_with_bundle_1_io_in_pre_decoder_jump),
    .io_in_pre_decoder_branchdata(Look_up_table_read_first_with_bundle_1_io_in_pre_decoder_branchdata),
    .io_in_pre_decoder_jr(Look_up_table_read_first_with_bundle_1_io_in_pre_decoder_jr),
    .io_in_true_branch_state(Look_up_table_read_first_with_bundle_1_io_in_true_branch_state),
    .io_out_pc(Look_up_table_read_first_with_bundle_1_io_out_pc),
    .io_out_inst(Look_up_table_read_first_with_bundle_1_io_out_inst),
    .io_out_exception_type(Look_up_table_read_first_with_bundle_1_io_out_exception_type),
    .io_out_pre_pc_target(Look_up_table_read_first_with_bundle_1_io_out_pre_pc_target),
    .io_out_pre_lookup_data(Look_up_table_read_first_with_bundle_1_io_out_pre_lookup_data),
    .io_out_pre_hashcode(Look_up_table_read_first_with_bundle_1_io_out_pre_hashcode),
    .io_out_pre_pht(Look_up_table_read_first_with_bundle_1_io_out_pre_pht),
    .io_out_pre_bht(Look_up_table_read_first_with_bundle_1_io_out_pre_bht),
    .io_out_pre_lookup_value(Look_up_table_read_first_with_bundle_1_io_out_pre_lookup_value),
    .io_out_pre_decoder_branchD_flag(Look_up_table_read_first_with_bundle_1_io_out_pre_decoder_branchD_flag),
    .io_out_pre_decoder_jump(Look_up_table_read_first_with_bundle_1_io_out_pre_decoder_jump),
    .io_out_pre_decoder_branchdata(Look_up_table_read_first_with_bundle_1_io_out_pre_decoder_branchdata),
    .io_out_pre_decoder_jr(Look_up_table_read_first_with_bundle_1_io_out_pre_decoder_jr),
    .io_out_true_branch_state(Look_up_table_read_first_with_bundle_1_io_out_true_branch_state)
  );
  Look_up_table_read_first_with_bundle Look_up_table_read_first_with_bundle_2 ( // @[fifo.scala 151:55]
    .clock(Look_up_table_read_first_with_bundle_2_clock),
    .reset(Look_up_table_read_first_with_bundle_2_reset),
    .io_ar_addr(Look_up_table_read_first_with_bundle_2_io_ar_addr),
    .io_aw_addr(Look_up_table_read_first_with_bundle_2_io_aw_addr),
    .io_write(Look_up_table_read_first_with_bundle_2_io_write),
    .io_in_pc(Look_up_table_read_first_with_bundle_2_io_in_pc),
    .io_in_inst(Look_up_table_read_first_with_bundle_2_io_in_inst),
    .io_in_pre_pc_target(Look_up_table_read_first_with_bundle_2_io_in_pre_pc_target),
    .io_in_pre_lookup_data(Look_up_table_read_first_with_bundle_2_io_in_pre_lookup_data),
    .io_in_pre_hashcode(Look_up_table_read_first_with_bundle_2_io_in_pre_hashcode),
    .io_in_pre_pht(Look_up_table_read_first_with_bundle_2_io_in_pre_pht),
    .io_in_pre_bht(Look_up_table_read_first_with_bundle_2_io_in_pre_bht),
    .io_in_pre_lookup_value(Look_up_table_read_first_with_bundle_2_io_in_pre_lookup_value),
    .io_in_pre_decoder_branchD_flag(Look_up_table_read_first_with_bundle_2_io_in_pre_decoder_branchD_flag),
    .io_in_pre_decoder_jump(Look_up_table_read_first_with_bundle_2_io_in_pre_decoder_jump),
    .io_in_pre_decoder_branchdata(Look_up_table_read_first_with_bundle_2_io_in_pre_decoder_branchdata),
    .io_in_pre_decoder_jr(Look_up_table_read_first_with_bundle_2_io_in_pre_decoder_jr),
    .io_in_true_branch_state(Look_up_table_read_first_with_bundle_2_io_in_true_branch_state),
    .io_out_pc(Look_up_table_read_first_with_bundle_2_io_out_pc),
    .io_out_inst(Look_up_table_read_first_with_bundle_2_io_out_inst),
    .io_out_exception_type(Look_up_table_read_first_with_bundle_2_io_out_exception_type),
    .io_out_pre_pc_target(Look_up_table_read_first_with_bundle_2_io_out_pre_pc_target),
    .io_out_pre_lookup_data(Look_up_table_read_first_with_bundle_2_io_out_pre_lookup_data),
    .io_out_pre_hashcode(Look_up_table_read_first_with_bundle_2_io_out_pre_hashcode),
    .io_out_pre_pht(Look_up_table_read_first_with_bundle_2_io_out_pre_pht),
    .io_out_pre_bht(Look_up_table_read_first_with_bundle_2_io_out_pre_bht),
    .io_out_pre_lookup_value(Look_up_table_read_first_with_bundle_2_io_out_pre_lookup_value),
    .io_out_pre_decoder_branchD_flag(Look_up_table_read_first_with_bundle_2_io_out_pre_decoder_branchD_flag),
    .io_out_pre_decoder_jump(Look_up_table_read_first_with_bundle_2_io_out_pre_decoder_jump),
    .io_out_pre_decoder_branchdata(Look_up_table_read_first_with_bundle_2_io_out_pre_decoder_branchdata),
    .io_out_pre_decoder_jr(Look_up_table_read_first_with_bundle_2_io_out_pre_decoder_jr),
    .io_out_true_branch_state(Look_up_table_read_first_with_bundle_2_io_out_true_branch_state)
  );
  Look_up_table_read_first_with_bundle Look_up_table_read_first_with_bundle_3 ( // @[fifo.scala 151:55]
    .clock(Look_up_table_read_first_with_bundle_3_clock),
    .reset(Look_up_table_read_first_with_bundle_3_reset),
    .io_ar_addr(Look_up_table_read_first_with_bundle_3_io_ar_addr),
    .io_aw_addr(Look_up_table_read_first_with_bundle_3_io_aw_addr),
    .io_write(Look_up_table_read_first_with_bundle_3_io_write),
    .io_in_pc(Look_up_table_read_first_with_bundle_3_io_in_pc),
    .io_in_inst(Look_up_table_read_first_with_bundle_3_io_in_inst),
    .io_in_pre_pc_target(Look_up_table_read_first_with_bundle_3_io_in_pre_pc_target),
    .io_in_pre_lookup_data(Look_up_table_read_first_with_bundle_3_io_in_pre_lookup_data),
    .io_in_pre_hashcode(Look_up_table_read_first_with_bundle_3_io_in_pre_hashcode),
    .io_in_pre_pht(Look_up_table_read_first_with_bundle_3_io_in_pre_pht),
    .io_in_pre_bht(Look_up_table_read_first_with_bundle_3_io_in_pre_bht),
    .io_in_pre_lookup_value(Look_up_table_read_first_with_bundle_3_io_in_pre_lookup_value),
    .io_in_pre_decoder_branchD_flag(Look_up_table_read_first_with_bundle_3_io_in_pre_decoder_branchD_flag),
    .io_in_pre_decoder_jump(Look_up_table_read_first_with_bundle_3_io_in_pre_decoder_jump),
    .io_in_pre_decoder_branchdata(Look_up_table_read_first_with_bundle_3_io_in_pre_decoder_branchdata),
    .io_in_pre_decoder_jr(Look_up_table_read_first_with_bundle_3_io_in_pre_decoder_jr),
    .io_in_true_branch_state(Look_up_table_read_first_with_bundle_3_io_in_true_branch_state),
    .io_out_pc(Look_up_table_read_first_with_bundle_3_io_out_pc),
    .io_out_inst(Look_up_table_read_first_with_bundle_3_io_out_inst),
    .io_out_exception_type(Look_up_table_read_first_with_bundle_3_io_out_exception_type),
    .io_out_pre_pc_target(Look_up_table_read_first_with_bundle_3_io_out_pre_pc_target),
    .io_out_pre_lookup_data(Look_up_table_read_first_with_bundle_3_io_out_pre_lookup_data),
    .io_out_pre_hashcode(Look_up_table_read_first_with_bundle_3_io_out_pre_hashcode),
    .io_out_pre_pht(Look_up_table_read_first_with_bundle_3_io_out_pre_pht),
    .io_out_pre_bht(Look_up_table_read_first_with_bundle_3_io_out_pre_bht),
    .io_out_pre_lookup_value(Look_up_table_read_first_with_bundle_3_io_out_pre_lookup_value),
    .io_out_pre_decoder_branchD_flag(Look_up_table_read_first_with_bundle_3_io_out_pre_decoder_branchD_flag),
    .io_out_pre_decoder_jump(Look_up_table_read_first_with_bundle_3_io_out_pre_decoder_jump),
    .io_out_pre_decoder_branchdata(Look_up_table_read_first_with_bundle_3_io_out_pre_decoder_branchdata),
    .io_out_pre_decoder_jr(Look_up_table_read_first_with_bundle_3_io_out_pre_decoder_jr),
    .io_out_true_branch_state(Look_up_table_read_first_with_bundle_3_io_out_true_branch_state)
  );
  assign io_read_out_0_pc = io_empty ? 64'h0 : _GEN_42; // @[fifo.scala 180:30]
  assign io_read_out_0_inst = io_empty ? 32'h0 : _GEN_43; // @[fifo.scala 180:30]
  assign io_read_out_0_exception_type = io_empty ? 2'h0 : _GEN_44; // @[fifo.scala 180:30]
  assign io_read_out_0_pre_pc_target = io_empty ? 64'h0 : _GEN_45; // @[fifo.scala 180:30]
  assign io_read_out_0_pre_lookup_data = io_empty ? 7'h0 : _GEN_46; // @[fifo.scala 180:30]
  assign io_read_out_0_pre_hashcode = io_empty ? 4'h0 : _GEN_47; // @[fifo.scala 180:30]
  assign io_read_out_0_pre_pht = io_empty ? 2'h0 : _GEN_48; // @[fifo.scala 180:30]
  assign io_read_out_0_pre_bht = io_empty ? 7'h0 : _GEN_49; // @[fifo.scala 180:30]
  assign io_read_out_0_pre_lookup_value = io_empty ? 8'h0 : _GEN_50; // @[fifo.scala 180:30]
  assign io_read_out_0_pre_decoder_branchD_flag = io_empty ? 1'h0 : _GEN_51; // @[fifo.scala 180:30]
  assign io_read_out_0_pre_decoder_jump = io_empty ? 1'h0 : _GEN_52; // @[fifo.scala 180:30]
  assign io_read_out_0_pre_decoder_branchdata = io_empty ? 6'h0 : _GEN_53; // @[fifo.scala 180:30]
  assign io_read_out_0_pre_decoder_jr = io_empty ? 1'h0 : _GEN_54; // @[fifo.scala 180:30]
  assign io_read_out_0_true_branch_state = io_empty ? 1'h0 : _GEN_55; // @[fifo.scala 180:30]
  assign io_full = _io_empty_T_1 ? _io_full_T_3 == _read_length_points_T_1 : _io_full_T_12; // @[fifo.scala 189:20]
  assign io_empty = write_banks_points == read_banks_points & write_length_points == read_length_points |
    io_point_write_en; // @[fifo.scala 187:106]
  assign Look_up_table_read_first_with_bundle_clock = clock;
  assign Look_up_table_read_first_with_bundle_reset = reset;
  assign Look_up_table_read_first_with_bundle_io_ar_addr = read_length_points; // @[fifo.scala 151:29 160:38]
  assign Look_up_table_read_first_with_bundle_io_aw_addr = write_length_points; // @[fifo.scala 151:29 159:38]
  assign Look_up_table_read_first_with_bundle_io_write = write_banks_points == 2'h0 & io_write_en[0]; // @[Mux.scala 81:58]
  assign Look_up_table_read_first_with_bundle_io_in_pc = io_write_in_0_pc; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_io_in_inst = io_write_in_0_inst; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_io_in_pre_pc_target = io_write_in_0_pre_pc_target; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_io_in_pre_lookup_data = io_write_in_0_pre_lookup_data; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_io_in_pre_hashcode = io_write_in_0_pre_hashcode; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_io_in_pre_pht = io_write_in_0_pre_pht; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_io_in_pre_bht = io_write_in_0_pre_bht; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_io_in_pre_lookup_value = io_write_in_0_pre_lookup_value; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_io_in_pre_decoder_branchD_flag = io_write_in_0_pre_decoder_branchD_flag; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_io_in_pre_decoder_jump = io_write_in_0_pre_decoder_jump; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_io_in_pre_decoder_branchdata = io_write_in_0_pre_decoder_branchdata; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_io_in_pre_decoder_jr = io_write_in_0_pre_decoder_jr; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_io_in_true_branch_state = io_write_in_0_true_branch_state; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_1_clock = clock;
  assign Look_up_table_read_first_with_bundle_1_reset = reset;
  assign Look_up_table_read_first_with_bundle_1_io_ar_addr = read_length_points; // @[fifo.scala 151:29 160:38]
  assign Look_up_table_read_first_with_bundle_1_io_aw_addr = write_length_points; // @[fifo.scala 151:29 159:38]
  assign Look_up_table_read_first_with_bundle_1_io_write = write_banks_points == 2'h1 & io_write_en[0]; // @[Mux.scala 81:58]
  assign Look_up_table_read_first_with_bundle_1_io_in_pc = io_write_in_0_pc; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_1_io_in_inst = io_write_in_0_inst; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_1_io_in_pre_pc_target = io_write_in_0_pre_pc_target; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_1_io_in_pre_lookup_data = io_write_in_0_pre_lookup_data; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_1_io_in_pre_hashcode = io_write_in_0_pre_hashcode; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_1_io_in_pre_pht = io_write_in_0_pre_pht; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_1_io_in_pre_bht = io_write_in_0_pre_bht; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_1_io_in_pre_lookup_value = io_write_in_0_pre_lookup_value; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_1_io_in_pre_decoder_branchD_flag = io_write_in_0_pre_decoder_branchD_flag; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_1_io_in_pre_decoder_jump = io_write_in_0_pre_decoder_jump; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_1_io_in_pre_decoder_branchdata = io_write_in_0_pre_decoder_branchdata; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_1_io_in_pre_decoder_jr = io_write_in_0_pre_decoder_jr; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_1_io_in_true_branch_state = io_write_in_0_true_branch_state; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_2_clock = clock;
  assign Look_up_table_read_first_with_bundle_2_reset = reset;
  assign Look_up_table_read_first_with_bundle_2_io_ar_addr = read_length_points; // @[fifo.scala 151:29 160:38]
  assign Look_up_table_read_first_with_bundle_2_io_aw_addr = write_length_points; // @[fifo.scala 151:29 159:38]
  assign Look_up_table_read_first_with_bundle_2_io_write = write_banks_points == 2'h2 & io_write_en[0]; // @[Mux.scala 81:58]
  assign Look_up_table_read_first_with_bundle_2_io_in_pc = io_write_in_0_pc; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_2_io_in_inst = io_write_in_0_inst; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_2_io_in_pre_pc_target = io_write_in_0_pre_pc_target; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_2_io_in_pre_lookup_data = io_write_in_0_pre_lookup_data; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_2_io_in_pre_hashcode = io_write_in_0_pre_hashcode; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_2_io_in_pre_pht = io_write_in_0_pre_pht; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_2_io_in_pre_bht = io_write_in_0_pre_bht; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_2_io_in_pre_lookup_value = io_write_in_0_pre_lookup_value; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_2_io_in_pre_decoder_branchD_flag = io_write_in_0_pre_decoder_branchD_flag; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_2_io_in_pre_decoder_jump = io_write_in_0_pre_decoder_jump; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_2_io_in_pre_decoder_branchdata = io_write_in_0_pre_decoder_branchdata; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_2_io_in_pre_decoder_jr = io_write_in_0_pre_decoder_jr; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_2_io_in_true_branch_state = io_write_in_0_true_branch_state; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_3_clock = clock;
  assign Look_up_table_read_first_with_bundle_3_reset = reset;
  assign Look_up_table_read_first_with_bundle_3_io_ar_addr = read_length_points; // @[fifo.scala 151:29 160:38]
  assign Look_up_table_read_first_with_bundle_3_io_aw_addr = write_length_points; // @[fifo.scala 151:29 159:38]
  assign Look_up_table_read_first_with_bundle_3_io_write = write_banks_points == 2'h3 & io_write_en[0]; // @[Mux.scala 81:58]
  assign Look_up_table_read_first_with_bundle_3_io_in_pc = io_write_in_0_pc; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_3_io_in_inst = io_write_in_0_inst; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_3_io_in_pre_pc_target = io_write_in_0_pre_pc_target; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_3_io_in_pre_lookup_data = io_write_in_0_pre_lookup_data; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_3_io_in_pre_hashcode = io_write_in_0_pre_hashcode; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_3_io_in_pre_pht = io_write_in_0_pre_pht; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_3_io_in_pre_bht = io_write_in_0_pre_bht; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_3_io_in_pre_lookup_value = io_write_in_0_pre_lookup_value; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_3_io_in_pre_decoder_branchD_flag = io_write_in_0_pre_decoder_branchD_flag; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_3_io_in_pre_decoder_jump = io_write_in_0_pre_decoder_jump; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_3_io_in_pre_decoder_branchdata = io_write_in_0_pre_decoder_branchdata; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_3_io_in_pre_decoder_jr = io_write_in_0_pre_decoder_jr; // @[fifo.scala 151:29 161:33]
  assign Look_up_table_read_first_with_bundle_3_io_in_true_branch_state = io_write_in_0_true_branch_state; // @[fifo.scala 151:29 161:33]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[fifo.scala 175:30]
      write_banks_points <= 2'h0;
    end else if (io_point_flush | io_point_write_en) begin
      write_banks_points <= 2'h0;
    end else begin
      write_banks_points <= _write_banks_points_T_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[fifo.scala 176:31]
      write_length_points <= 4'h0;
    end else if (_write_banks_points_T) begin
      write_length_points <= 4'h0;
    end else begin
      write_length_points <= _write_length_points_T_7;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[fifo.scala 177:29]
      read_banks_points <= 2'h0;
    end else if (_write_banks_points_T) begin
      read_banks_points <= 2'h0;
    end else begin
      read_banks_points <= _read_banks_points_T_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[fifo.scala 178:30]
      read_length_points <= 4'h0;
    end else if (_write_banks_points_T) begin
      read_length_points <= 4'h0;
    end else begin
      read_length_points <= _read_length_points_T_7;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  write_banks_points = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  write_length_points = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  read_banks_points = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  read_length_points = _RAND_3[3:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    write_banks_points = 2'h0;
  end
  if (reset) begin
    write_length_points = 4'h0;
  end
  if (reset) begin
    read_banks_points = 2'h0;
  end
  if (reset) begin
    read_length_points = 4'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module pc_detail(
  input         clock,
  input         reset,
  input         io_stall,
  input         io_flush,
  input  [63:0] io_in_pc_value_in,
  output [63:0] io_out_pc_value_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] pc_value; // @[myCPU.scala 325:25]
  assign io_out_pc_value_out = pc_value; // @[myCPU.scala 328:25]
  always @(posedge clock) begin
    if (reset) begin // @[myCPU.scala 327:20]
      pc_value <= 64'h7ffffffc;
    end else if (io_flush) begin // @[myCPU.scala 327:60]
      pc_value <= 64'h0;
    end else if (io_stall) begin // @[myCPU.scala 327:77]
      pc_value <= io_in_pc_value_in;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc_value = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Look_up_table_read_first_(
  input        clock,
  input        reset,
  input  [4:0] io_ar_addr,
  input  [4:0] io_aw_addr,
  input        io_write,
  input  [7:0] io_in,
  output [7:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] btb_0; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_1; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_2; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_3; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_4; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_5; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_6; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_7; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_8; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_9; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_10; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_11; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_12; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_13; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_14; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_15; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_16; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_17; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_18; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_19; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_20; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_21; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_22; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_23; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_24; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_25; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_26; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_27; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_28; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_29; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_30; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_31; // @[ports_lookup_table.scala 81:22]
  wire [7:0] _GEN_1 = 5'h1 == io_ar_addr ? btb_1 : btb_0; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_2 = 5'h2 == io_ar_addr ? btb_2 : _GEN_1; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_3 = 5'h3 == io_ar_addr ? btb_3 : _GEN_2; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_4 = 5'h4 == io_ar_addr ? btb_4 : _GEN_3; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_5 = 5'h5 == io_ar_addr ? btb_5 : _GEN_4; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_6 = 5'h6 == io_ar_addr ? btb_6 : _GEN_5; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_7 = 5'h7 == io_ar_addr ? btb_7 : _GEN_6; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_8 = 5'h8 == io_ar_addr ? btb_8 : _GEN_7; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_9 = 5'h9 == io_ar_addr ? btb_9 : _GEN_8; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_10 = 5'ha == io_ar_addr ? btb_10 : _GEN_9; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_11 = 5'hb == io_ar_addr ? btb_11 : _GEN_10; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_12 = 5'hc == io_ar_addr ? btb_12 : _GEN_11; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_13 = 5'hd == io_ar_addr ? btb_13 : _GEN_12; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_14 = 5'he == io_ar_addr ? btb_14 : _GEN_13; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_15 = 5'hf == io_ar_addr ? btb_15 : _GEN_14; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_16 = 5'h10 == io_ar_addr ? btb_16 : _GEN_15; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_17 = 5'h11 == io_ar_addr ? btb_17 : _GEN_16; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_18 = 5'h12 == io_ar_addr ? btb_18 : _GEN_17; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_19 = 5'h13 == io_ar_addr ? btb_19 : _GEN_18; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_20 = 5'h14 == io_ar_addr ? btb_20 : _GEN_19; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_21 = 5'h15 == io_ar_addr ? btb_21 : _GEN_20; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_22 = 5'h16 == io_ar_addr ? btb_22 : _GEN_21; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_23 = 5'h17 == io_ar_addr ? btb_23 : _GEN_22; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_24 = 5'h18 == io_ar_addr ? btb_24 : _GEN_23; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_25 = 5'h19 == io_ar_addr ? btb_25 : _GEN_24; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_26 = 5'h1a == io_ar_addr ? btb_26 : _GEN_25; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_27 = 5'h1b == io_ar_addr ? btb_27 : _GEN_26; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_28 = 5'h1c == io_ar_addr ? btb_28 : _GEN_27; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_29 = 5'h1d == io_ar_addr ? btb_29 : _GEN_28; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_30 = 5'h1e == io_ar_addr ? btb_30 : _GEN_29; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_33 = 5'h1 == io_aw_addr ? btb_1 : btb_0; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_34 = 5'h2 == io_aw_addr ? btb_2 : _GEN_33; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_35 = 5'h3 == io_aw_addr ? btb_3 : _GEN_34; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_36 = 5'h4 == io_aw_addr ? btb_4 : _GEN_35; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_37 = 5'h5 == io_aw_addr ? btb_5 : _GEN_36; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_38 = 5'h6 == io_aw_addr ? btb_6 : _GEN_37; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_39 = 5'h7 == io_aw_addr ? btb_7 : _GEN_38; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_40 = 5'h8 == io_aw_addr ? btb_8 : _GEN_39; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_41 = 5'h9 == io_aw_addr ? btb_9 : _GEN_40; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_42 = 5'ha == io_aw_addr ? btb_10 : _GEN_41; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_43 = 5'hb == io_aw_addr ? btb_11 : _GEN_42; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_44 = 5'hc == io_aw_addr ? btb_12 : _GEN_43; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_45 = 5'hd == io_aw_addr ? btb_13 : _GEN_44; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_46 = 5'he == io_aw_addr ? btb_14 : _GEN_45; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_47 = 5'hf == io_aw_addr ? btb_15 : _GEN_46; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_48 = 5'h10 == io_aw_addr ? btb_16 : _GEN_47; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_49 = 5'h11 == io_aw_addr ? btb_17 : _GEN_48; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_50 = 5'h12 == io_aw_addr ? btb_18 : _GEN_49; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_51 = 5'h13 == io_aw_addr ? btb_19 : _GEN_50; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_52 = 5'h14 == io_aw_addr ? btb_20 : _GEN_51; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_53 = 5'h15 == io_aw_addr ? btb_21 : _GEN_52; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_54 = 5'h16 == io_aw_addr ? btb_22 : _GEN_53; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_55 = 5'h17 == io_aw_addr ? btb_23 : _GEN_54; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_56 = 5'h18 == io_aw_addr ? btb_24 : _GEN_55; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_57 = 5'h19 == io_aw_addr ? btb_25 : _GEN_56; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_58 = 5'h1a == io_aw_addr ? btb_26 : _GEN_57; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_59 = 5'h1b == io_aw_addr ? btb_27 : _GEN_58; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_60 = 5'h1c == io_aw_addr ? btb_28 : _GEN_59; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_61 = 5'h1d == io_aw_addr ? btb_29 : _GEN_60; // @[ports_lookup_table.scala 83:{27,27}]
  assign io_out = 5'h1f == io_ar_addr ? btb_31 : _GEN_30; // @[ports_lookup_table.scala 82:{12,12}]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_0 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_0 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_0 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_0 <= btb_30;
      end else begin
        btb_0 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_1 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_1 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_1 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_1 <= btb_30;
      end else begin
        btb_1 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_2 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_2 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_2 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_2 <= btb_30;
      end else begin
        btb_2 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_3 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_3 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_3 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_3 <= btb_30;
      end else begin
        btb_3 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_4 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_4 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_4 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_4 <= btb_30;
      end else begin
        btb_4 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_5 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_5 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_5 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_5 <= btb_30;
      end else begin
        btb_5 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_6 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_6 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_6 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_6 <= btb_30;
      end else begin
        btb_6 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_7 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_7 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_7 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_7 <= btb_30;
      end else begin
        btb_7 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_8 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_8 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_8 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_8 <= btb_30;
      end else begin
        btb_8 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_9 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_9 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_9 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_9 <= btb_30;
      end else begin
        btb_9 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_10 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'ha == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_10 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_10 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_10 <= btb_30;
      end else begin
        btb_10 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_11 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'hb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_11 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_11 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_11 <= btb_30;
      end else begin
        btb_11 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_12 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'hc == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_12 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_12 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_12 <= btb_30;
      end else begin
        btb_12 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_13 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'hd == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_13 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_13 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_13 <= btb_30;
      end else begin
        btb_13 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_14 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'he == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_14 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_14 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_14 <= btb_30;
      end else begin
        btb_14 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_15 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'hf == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_15 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_15 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_15 <= btb_30;
      end else begin
        btb_15 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_16 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h10 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_16 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_16 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_16 <= btb_30;
      end else begin
        btb_16 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_17 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h11 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_17 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_17 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_17 <= btb_30;
      end else begin
        btb_17 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_18 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h12 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_18 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_18 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_18 <= btb_30;
      end else begin
        btb_18 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_19 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h13 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_19 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_19 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_19 <= btb_30;
      end else begin
        btb_19 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_20 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h14 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_20 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_20 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_20 <= btb_30;
      end else begin
        btb_20 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_21 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h15 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_21 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_21 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_21 <= btb_30;
      end else begin
        btb_21 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_22 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h16 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_22 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_22 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_22 <= btb_30;
      end else begin
        btb_22 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_23 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h17 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_23 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_23 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_23 <= btb_30;
      end else begin
        btb_23 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_24 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h18 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_24 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_24 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_24 <= btb_30;
      end else begin
        btb_24 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_25 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h19 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_25 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_25 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_25 <= btb_30;
      end else begin
        btb_25 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_26 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h1a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_26 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_26 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_26 <= btb_30;
      end else begin
        btb_26 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_27 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h1b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_27 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_27 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_27 <= btb_30;
      end else begin
        btb_27 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_28 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h1c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_28 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_28 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_28 <= btb_30;
      end else begin
        btb_28 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_29 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h1d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_29 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_29 <= btb_31;
      end else if (5'h1e == io_aw_addr) begin
        btb_29 <= btb_30;
      end else begin
        btb_29 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_30 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h1e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_30 <= io_in;
      end else if (5'h1f == io_aw_addr) begin
        btb_30 <= btb_31;
      end else if (!(5'h1e == io_aw_addr)) begin
        btb_30 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_31 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (5'h1f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_31 <= io_in;
      end else if (!(5'h1f == io_aw_addr)) begin
        if (5'h1e == io_aw_addr) begin
          btb_31 <= btb_30;
        end else begin
          btb_31 <= _GEN_61;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  btb_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  btb_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  btb_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  btb_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  btb_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  btb_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  btb_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  btb_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  btb_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  btb_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  btb_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  btb_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  btb_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  btb_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  btb_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  btb_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  btb_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  btb_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  btb_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  btb_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  btb_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  btb_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  btb_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  btb_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  btb_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  btb_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  btb_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  btb_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  btb_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  btb_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  btb_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  btb_31 = _RAND_31[7:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    btb_0 = 8'h0;
  end
  if (reset) begin
    btb_1 = 8'h0;
  end
  if (reset) begin
    btb_2 = 8'h0;
  end
  if (reset) begin
    btb_3 = 8'h0;
  end
  if (reset) begin
    btb_4 = 8'h0;
  end
  if (reset) begin
    btb_5 = 8'h0;
  end
  if (reset) begin
    btb_6 = 8'h0;
  end
  if (reset) begin
    btb_7 = 8'h0;
  end
  if (reset) begin
    btb_8 = 8'h0;
  end
  if (reset) begin
    btb_9 = 8'h0;
  end
  if (reset) begin
    btb_10 = 8'h0;
  end
  if (reset) begin
    btb_11 = 8'h0;
  end
  if (reset) begin
    btb_12 = 8'h0;
  end
  if (reset) begin
    btb_13 = 8'h0;
  end
  if (reset) begin
    btb_14 = 8'h0;
  end
  if (reset) begin
    btb_15 = 8'h0;
  end
  if (reset) begin
    btb_16 = 8'h0;
  end
  if (reset) begin
    btb_17 = 8'h0;
  end
  if (reset) begin
    btb_18 = 8'h0;
  end
  if (reset) begin
    btb_19 = 8'h0;
  end
  if (reset) begin
    btb_20 = 8'h0;
  end
  if (reset) begin
    btb_21 = 8'h0;
  end
  if (reset) begin
    btb_22 = 8'h0;
  end
  if (reset) begin
    btb_23 = 8'h0;
  end
  if (reset) begin
    btb_24 = 8'h0;
  end
  if (reset) begin
    btb_25 = 8'h0;
  end
  if (reset) begin
    btb_26 = 8'h0;
  end
  if (reset) begin
    btb_27 = 8'h0;
  end
  if (reset) begin
    btb_28 = 8'h0;
  end
  if (reset) begin
    btb_29 = 8'h0;
  end
  if (reset) begin
    btb_30 = 8'h0;
  end
  if (reset) begin
    btb_31 = 8'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module data_ram_simple_two_ports(
  input        clock,
  input        reset,
  input        io_wea,
  input  [4:0] io_addra,
  input  [7:0] io_dina,
  input  [4:0] io_addrb,
  output [7:0] io_doutb
);
  wire  Look_up_table_read_first__clock; // @[ip_user.scala 97:23]
  wire  Look_up_table_read_first__reset; // @[ip_user.scala 97:23]
  wire [4:0] Look_up_table_read_first__io_ar_addr; // @[ip_user.scala 97:23]
  wire [4:0] Look_up_table_read_first__io_aw_addr; // @[ip_user.scala 97:23]
  wire  Look_up_table_read_first__io_write; // @[ip_user.scala 97:23]
  wire [7:0] Look_up_table_read_first__io_in; // @[ip_user.scala 97:23]
  wire [7:0] Look_up_table_read_first__io_out; // @[ip_user.scala 97:23]
  Look_up_table_read_first_ Look_up_table_read_first_ ( // @[ip_user.scala 97:23]
    .clock(Look_up_table_read_first__clock),
    .reset(Look_up_table_read_first__reset),
    .io_ar_addr(Look_up_table_read_first__io_ar_addr),
    .io_aw_addr(Look_up_table_read_first__io_aw_addr),
    .io_write(Look_up_table_read_first__io_write),
    .io_in(Look_up_table_read_first__io_in),
    .io_out(Look_up_table_read_first__io_out)
  );
  assign io_doutb = Look_up_table_read_first__io_out; // @[ip_user.scala 102:19]
  assign Look_up_table_read_first__clock = clock;
  assign Look_up_table_read_first__reset = reset;
  assign Look_up_table_read_first__io_ar_addr = io_addra; // @[ip_user.scala 98:19]
  assign Look_up_table_read_first__io_aw_addr = io_addrb; // @[ip_user.scala 99:19]
  assign Look_up_table_read_first__io_write = io_wea; // @[ip_user.scala 101:19]
  assign Look_up_table_read_first__io_in = io_dina; // @[ip_user.scala 100:19]
endmodule
module pht_data_with_block_ram(
  input        clock,
  input        reset,
  input        io_wen,
  input  [4:0] io_raddr,
  input  [4:0] io_waddr,
  input  [7:0] io_wdata,
  output [7:0] io_rdata
);
  wire  btb_data_ram_0_clock; // @[PHTS.scala 176:32]
  wire  btb_data_ram_0_reset; // @[PHTS.scala 176:32]
  wire  btb_data_ram_0_io_wea; // @[PHTS.scala 176:32]
  wire [4:0] btb_data_ram_0_io_addra; // @[PHTS.scala 176:32]
  wire [7:0] btb_data_ram_0_io_dina; // @[PHTS.scala 176:32]
  wire [4:0] btb_data_ram_0_io_addrb; // @[PHTS.scala 176:32]
  wire [7:0] btb_data_ram_0_io_doutb; // @[PHTS.scala 176:32]
  data_ram_simple_two_ports btb_data_ram_0 ( // @[PHTS.scala 176:32]
    .clock(btb_data_ram_0_clock),
    .reset(btb_data_ram_0_reset),
    .io_wea(btb_data_ram_0_io_wea),
    .io_addra(btb_data_ram_0_io_addra),
    .io_dina(btb_data_ram_0_io_dina),
    .io_addrb(btb_data_ram_0_io_addrb),
    .io_doutb(btb_data_ram_0_io_doutb)
  );
  assign io_rdata = btb_data_ram_0_io_doutb; // @[PHTS.scala 185:18]
  assign btb_data_ram_0_clock = clock;
  assign btb_data_ram_0_reset = reset;
  assign btb_data_ram_0_io_wea = io_wen; // @[PHTS.scala 181:28]
  assign btb_data_ram_0_io_addra = io_waddr; // @[PHTS.scala 182:29]
  assign btb_data_ram_0_io_dina = io_wdata; // @[PHTS.scala 184:28]
  assign btb_data_ram_0_io_addrb = io_raddr; // @[PHTS.scala 183:29]
endmodule
module PHTS_with_block_ram(
  input        clock,
  input        reset,
  input  [6:0] io_ar_addr,
  input  [2:0] io_ar_pht_addr,
  input  [6:0] io_aw_addr,
  input  [2:0] io_aw_pht_addr,
  input        io_write,
  input  [7:0] io_in,
  output [7:0] io_pht_out,
  output [1:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  pht_data_with_block_ram_clock; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_reset; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_io_wen; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_io_raddr; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_io_waddr; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_io_wdata; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_io_rdata; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_1_clock; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_1_reset; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_1_io_wen; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_1_io_raddr; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_1_io_waddr; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_1_io_wdata; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_1_io_rdata; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_2_clock; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_2_reset; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_2_io_wen; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_2_io_raddr; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_2_io_waddr; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_2_io_wdata; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_2_io_rdata; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_3_clock; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_3_reset; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_3_io_wen; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_3_io_raddr; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_3_io_waddr; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_3_io_wdata; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_3_io_rdata; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_4_clock; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_4_reset; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_4_io_wen; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_4_io_raddr; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_4_io_waddr; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_4_io_wdata; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_4_io_rdata; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_5_clock; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_5_reset; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_5_io_wen; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_5_io_raddr; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_5_io_waddr; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_5_io_wdata; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_5_io_rdata; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_6_clock; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_6_reset; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_6_io_wen; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_6_io_raddr; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_6_io_waddr; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_6_io_wdata; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_6_io_rdata; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_7_clock; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_7_reset; // @[PHTS.scala 205:45]
  wire  pht_data_with_block_ram_7_io_wen; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_7_io_raddr; // @[PHTS.scala 205:45]
  wire [4:0] pht_data_with_block_ram_7_io_waddr; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_7_io_wdata; // @[PHTS.scala 205:45]
  wire [7:0] pht_data_with_block_ram_7_io_rdata; // @[PHTS.scala 205:45]
  reg [6:0] raddr_reg; // @[PHTS.scala 213:28]
  reg [7:0] ways_araddr_reg; // @[PHTS.scala 214:34]
  wire [7:0] phts_0_rdata = pht_data_with_block_ram_io_rdata; // @[PHTS.scala 205:{23,23}]
  wire [7:0] phts_1_rdata = pht_data_with_block_ram_1_io_rdata; // @[PHTS.scala 205:{23,23}]
  wire [7:0] _GEN_1 = 3'h1 == ways_araddr_reg[2:0] ? phts_1_rdata : phts_0_rdata; // @[PHTS.scala 217:{67,67}]
  wire [7:0] phts_2_rdata = pht_data_with_block_ram_2_io_rdata; // @[PHTS.scala 205:{23,23}]
  wire [7:0] _GEN_2 = 3'h2 == ways_araddr_reg[2:0] ? phts_2_rdata : _GEN_1; // @[PHTS.scala 217:{67,67}]
  wire [7:0] phts_3_rdata = pht_data_with_block_ram_3_io_rdata; // @[PHTS.scala 205:{23,23}]
  wire [7:0] _GEN_3 = 3'h3 == ways_araddr_reg[2:0] ? phts_3_rdata : _GEN_2; // @[PHTS.scala 217:{67,67}]
  wire [7:0] phts_4_rdata = pht_data_with_block_ram_4_io_rdata; // @[PHTS.scala 205:{23,23}]
  wire [7:0] _GEN_4 = 3'h4 == ways_araddr_reg[2:0] ? phts_4_rdata : _GEN_3; // @[PHTS.scala 217:{67,67}]
  wire [7:0] phts_5_rdata = pht_data_with_block_ram_5_io_rdata; // @[PHTS.scala 205:{23,23}]
  wire [7:0] _GEN_5 = 3'h5 == ways_araddr_reg[2:0] ? phts_5_rdata : _GEN_4; // @[PHTS.scala 217:{67,67}]
  wire [7:0] phts_6_rdata = pht_data_with_block_ram_6_io_rdata; // @[PHTS.scala 205:{23,23}]
  wire [7:0] _GEN_6 = 3'h6 == ways_araddr_reg[2:0] ? phts_6_rdata : _GEN_5; // @[PHTS.scala 217:{67,67}]
  wire [7:0] phts_7_rdata = pht_data_with_block_ram_7_io_rdata; // @[PHTS.scala 205:{23,23}]
  wire [7:0] _GEN_7 = 3'h7 == ways_araddr_reg[2:0] ? phts_7_rdata : _GEN_6; // @[PHTS.scala 217:{67,67}]
  wire [1:0] _io_out_T_10 = 2'h0 == raddr_reg[1:0] ? _GEN_7[1:0] : _GEN_7[7:6]; // @[Mux.scala 81:58]
  wire [1:0] _io_out_T_12 = 2'h1 == raddr_reg[1:0] ? _GEN_7[3:2] : _io_out_T_10; // @[Mux.scala 81:58]
  pht_data_with_block_ram pht_data_with_block_ram ( // @[PHTS.scala 205:45]
    .clock(pht_data_with_block_ram_clock),
    .reset(pht_data_with_block_ram_reset),
    .io_wen(pht_data_with_block_ram_io_wen),
    .io_raddr(pht_data_with_block_ram_io_raddr),
    .io_waddr(pht_data_with_block_ram_io_waddr),
    .io_wdata(pht_data_with_block_ram_io_wdata),
    .io_rdata(pht_data_with_block_ram_io_rdata)
  );
  pht_data_with_block_ram pht_data_with_block_ram_1 ( // @[PHTS.scala 205:45]
    .clock(pht_data_with_block_ram_1_clock),
    .reset(pht_data_with_block_ram_1_reset),
    .io_wen(pht_data_with_block_ram_1_io_wen),
    .io_raddr(pht_data_with_block_ram_1_io_raddr),
    .io_waddr(pht_data_with_block_ram_1_io_waddr),
    .io_wdata(pht_data_with_block_ram_1_io_wdata),
    .io_rdata(pht_data_with_block_ram_1_io_rdata)
  );
  pht_data_with_block_ram pht_data_with_block_ram_2 ( // @[PHTS.scala 205:45]
    .clock(pht_data_with_block_ram_2_clock),
    .reset(pht_data_with_block_ram_2_reset),
    .io_wen(pht_data_with_block_ram_2_io_wen),
    .io_raddr(pht_data_with_block_ram_2_io_raddr),
    .io_waddr(pht_data_with_block_ram_2_io_waddr),
    .io_wdata(pht_data_with_block_ram_2_io_wdata),
    .io_rdata(pht_data_with_block_ram_2_io_rdata)
  );
  pht_data_with_block_ram pht_data_with_block_ram_3 ( // @[PHTS.scala 205:45]
    .clock(pht_data_with_block_ram_3_clock),
    .reset(pht_data_with_block_ram_3_reset),
    .io_wen(pht_data_with_block_ram_3_io_wen),
    .io_raddr(pht_data_with_block_ram_3_io_raddr),
    .io_waddr(pht_data_with_block_ram_3_io_waddr),
    .io_wdata(pht_data_with_block_ram_3_io_wdata),
    .io_rdata(pht_data_with_block_ram_3_io_rdata)
  );
  pht_data_with_block_ram pht_data_with_block_ram_4 ( // @[PHTS.scala 205:45]
    .clock(pht_data_with_block_ram_4_clock),
    .reset(pht_data_with_block_ram_4_reset),
    .io_wen(pht_data_with_block_ram_4_io_wen),
    .io_raddr(pht_data_with_block_ram_4_io_raddr),
    .io_waddr(pht_data_with_block_ram_4_io_waddr),
    .io_wdata(pht_data_with_block_ram_4_io_wdata),
    .io_rdata(pht_data_with_block_ram_4_io_rdata)
  );
  pht_data_with_block_ram pht_data_with_block_ram_5 ( // @[PHTS.scala 205:45]
    .clock(pht_data_with_block_ram_5_clock),
    .reset(pht_data_with_block_ram_5_reset),
    .io_wen(pht_data_with_block_ram_5_io_wen),
    .io_raddr(pht_data_with_block_ram_5_io_raddr),
    .io_waddr(pht_data_with_block_ram_5_io_waddr),
    .io_wdata(pht_data_with_block_ram_5_io_wdata),
    .io_rdata(pht_data_with_block_ram_5_io_rdata)
  );
  pht_data_with_block_ram pht_data_with_block_ram_6 ( // @[PHTS.scala 205:45]
    .clock(pht_data_with_block_ram_6_clock),
    .reset(pht_data_with_block_ram_6_reset),
    .io_wen(pht_data_with_block_ram_6_io_wen),
    .io_raddr(pht_data_with_block_ram_6_io_raddr),
    .io_waddr(pht_data_with_block_ram_6_io_waddr),
    .io_wdata(pht_data_with_block_ram_6_io_wdata),
    .io_rdata(pht_data_with_block_ram_6_io_rdata)
  );
  pht_data_with_block_ram pht_data_with_block_ram_7 ( // @[PHTS.scala 205:45]
    .clock(pht_data_with_block_ram_7_clock),
    .reset(pht_data_with_block_ram_7_reset),
    .io_wen(pht_data_with_block_ram_7_io_wen),
    .io_raddr(pht_data_with_block_ram_7_io_raddr),
    .io_waddr(pht_data_with_block_ram_7_io_waddr),
    .io_wdata(pht_data_with_block_ram_7_io_wdata),
    .io_rdata(pht_data_with_block_ram_7_io_rdata)
  );
  assign io_pht_out = 3'h7 == ways_araddr_reg[2:0] ? phts_7_rdata : _GEN_6; // @[PHTS.scala 222:{16,16}]
  assign io_out = 2'h2 == raddr_reg[1:0] ? _GEN_7[5:4] : _io_out_T_12; // @[Mux.scala 81:58]
  assign pht_data_with_block_ram_clock = clock;
  assign pht_data_with_block_ram_reset = reset;
  assign pht_data_with_block_ram_io_wen = io_aw_pht_addr == 3'h0 & io_write; // @[PHTS.scala 207:52]
  assign pht_data_with_block_ram_io_raddr = io_ar_addr[6:2]; // @[PHTS.scala 210:36]
  assign pht_data_with_block_ram_io_waddr = io_aw_addr[6:2]; // @[PHTS.scala 211:36]
  assign pht_data_with_block_ram_io_wdata = io_in; // @[PHTS.scala 205:23 209:23]
  assign pht_data_with_block_ram_1_clock = clock;
  assign pht_data_with_block_ram_1_reset = reset;
  assign pht_data_with_block_ram_1_io_wen = io_aw_pht_addr == 3'h1 & io_write; // @[PHTS.scala 207:52]
  assign pht_data_with_block_ram_1_io_raddr = io_ar_addr[6:2]; // @[PHTS.scala 210:36]
  assign pht_data_with_block_ram_1_io_waddr = io_aw_addr[6:2]; // @[PHTS.scala 211:36]
  assign pht_data_with_block_ram_1_io_wdata = io_in; // @[PHTS.scala 205:23 209:23]
  assign pht_data_with_block_ram_2_clock = clock;
  assign pht_data_with_block_ram_2_reset = reset;
  assign pht_data_with_block_ram_2_io_wen = io_aw_pht_addr == 3'h2 & io_write; // @[PHTS.scala 207:52]
  assign pht_data_with_block_ram_2_io_raddr = io_ar_addr[6:2]; // @[PHTS.scala 210:36]
  assign pht_data_with_block_ram_2_io_waddr = io_aw_addr[6:2]; // @[PHTS.scala 211:36]
  assign pht_data_with_block_ram_2_io_wdata = io_in; // @[PHTS.scala 205:23 209:23]
  assign pht_data_with_block_ram_3_clock = clock;
  assign pht_data_with_block_ram_3_reset = reset;
  assign pht_data_with_block_ram_3_io_wen = io_aw_pht_addr == 3'h3 & io_write; // @[PHTS.scala 207:52]
  assign pht_data_with_block_ram_3_io_raddr = io_ar_addr[6:2]; // @[PHTS.scala 210:36]
  assign pht_data_with_block_ram_3_io_waddr = io_aw_addr[6:2]; // @[PHTS.scala 211:36]
  assign pht_data_with_block_ram_3_io_wdata = io_in; // @[PHTS.scala 205:23 209:23]
  assign pht_data_with_block_ram_4_clock = clock;
  assign pht_data_with_block_ram_4_reset = reset;
  assign pht_data_with_block_ram_4_io_wen = io_aw_pht_addr == 3'h4 & io_write; // @[PHTS.scala 207:52]
  assign pht_data_with_block_ram_4_io_raddr = io_ar_addr[6:2]; // @[PHTS.scala 210:36]
  assign pht_data_with_block_ram_4_io_waddr = io_aw_addr[6:2]; // @[PHTS.scala 211:36]
  assign pht_data_with_block_ram_4_io_wdata = io_in; // @[PHTS.scala 205:23 209:23]
  assign pht_data_with_block_ram_5_clock = clock;
  assign pht_data_with_block_ram_5_reset = reset;
  assign pht_data_with_block_ram_5_io_wen = io_aw_pht_addr == 3'h5 & io_write; // @[PHTS.scala 207:52]
  assign pht_data_with_block_ram_5_io_raddr = io_ar_addr[6:2]; // @[PHTS.scala 210:36]
  assign pht_data_with_block_ram_5_io_waddr = io_aw_addr[6:2]; // @[PHTS.scala 211:36]
  assign pht_data_with_block_ram_5_io_wdata = io_in; // @[PHTS.scala 205:23 209:23]
  assign pht_data_with_block_ram_6_clock = clock;
  assign pht_data_with_block_ram_6_reset = reset;
  assign pht_data_with_block_ram_6_io_wen = io_aw_pht_addr == 3'h6 & io_write; // @[PHTS.scala 207:52]
  assign pht_data_with_block_ram_6_io_raddr = io_ar_addr[6:2]; // @[PHTS.scala 210:36]
  assign pht_data_with_block_ram_6_io_waddr = io_aw_addr[6:2]; // @[PHTS.scala 211:36]
  assign pht_data_with_block_ram_6_io_wdata = io_in; // @[PHTS.scala 205:23 209:23]
  assign pht_data_with_block_ram_7_clock = clock;
  assign pht_data_with_block_ram_7_reset = reset;
  assign pht_data_with_block_ram_7_io_wen = io_aw_pht_addr == 3'h7 & io_write; // @[PHTS.scala 207:52]
  assign pht_data_with_block_ram_7_io_raddr = io_ar_addr[6:2]; // @[PHTS.scala 210:36]
  assign pht_data_with_block_ram_7_io_waddr = io_aw_addr[6:2]; // @[PHTS.scala 211:36]
  assign pht_data_with_block_ram_7_io_wdata = io_in; // @[PHTS.scala 205:23 209:23]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PHTS.scala 213:28]
      raddr_reg <= 7'h0; // @[PHTS.scala 213:28]
    end else begin
      raddr_reg <= io_ar_addr; // @[PHTS.scala 215:15]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PHTS.scala 214:34]
      ways_araddr_reg <= 8'h0; // @[PHTS.scala 214:34]
    end else begin
      ways_araddr_reg <= {{5'd0}, io_ar_pht_addr}; // @[PHTS.scala 216:21]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  raddr_reg = _RAND_0[6:0];
  _RAND_1 = {1{`RANDOM}};
  ways_araddr_reg = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    raddr_reg = 7'h0;
  end
  if (reset) begin
    ways_araddr_reg = 8'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PHTS_banks_oneissue_block_ram(
  input        clock,
  input        reset,
  input  [1:0] io_ar_bank_sel,
  input  [6:0] io_ar_addr_L,
  input  [2:0] io_ar_pht_addr,
  input  [6:0] io_aw_addr,
  input  [2:0] io_aw_pht_addr,
  input  [1:0] io_aw_bank_sel,
  input        io_write,
  input  [7:0] io_in,
  output [1:0] io_out_L,
  output [7:0] io_pht_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  PHTS_with_block_ram_clock; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_reset; // @[PHTS.scala 250:55]
  wire [6:0] PHTS_with_block_ram_io_ar_addr; // @[PHTS.scala 250:55]
  wire [2:0] PHTS_with_block_ram_io_ar_pht_addr; // @[PHTS.scala 250:55]
  wire [6:0] PHTS_with_block_ram_io_aw_addr; // @[PHTS.scala 250:55]
  wire [2:0] PHTS_with_block_ram_io_aw_pht_addr; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_io_write; // @[PHTS.scala 250:55]
  wire [7:0] PHTS_with_block_ram_io_in; // @[PHTS.scala 250:55]
  wire [7:0] PHTS_with_block_ram_io_pht_out; // @[PHTS.scala 250:55]
  wire [1:0] PHTS_with_block_ram_io_out; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_1_clock; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_1_reset; // @[PHTS.scala 250:55]
  wire [6:0] PHTS_with_block_ram_1_io_ar_addr; // @[PHTS.scala 250:55]
  wire [2:0] PHTS_with_block_ram_1_io_ar_pht_addr; // @[PHTS.scala 250:55]
  wire [6:0] PHTS_with_block_ram_1_io_aw_addr; // @[PHTS.scala 250:55]
  wire [2:0] PHTS_with_block_ram_1_io_aw_pht_addr; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_1_io_write; // @[PHTS.scala 250:55]
  wire [7:0] PHTS_with_block_ram_1_io_in; // @[PHTS.scala 250:55]
  wire [7:0] PHTS_with_block_ram_1_io_pht_out; // @[PHTS.scala 250:55]
  wire [1:0] PHTS_with_block_ram_1_io_out; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_2_clock; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_2_reset; // @[PHTS.scala 250:55]
  wire [6:0] PHTS_with_block_ram_2_io_ar_addr; // @[PHTS.scala 250:55]
  wire [2:0] PHTS_with_block_ram_2_io_ar_pht_addr; // @[PHTS.scala 250:55]
  wire [6:0] PHTS_with_block_ram_2_io_aw_addr; // @[PHTS.scala 250:55]
  wire [2:0] PHTS_with_block_ram_2_io_aw_pht_addr; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_2_io_write; // @[PHTS.scala 250:55]
  wire [7:0] PHTS_with_block_ram_2_io_in; // @[PHTS.scala 250:55]
  wire [7:0] PHTS_with_block_ram_2_io_pht_out; // @[PHTS.scala 250:55]
  wire [1:0] PHTS_with_block_ram_2_io_out; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_3_clock; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_3_reset; // @[PHTS.scala 250:55]
  wire [6:0] PHTS_with_block_ram_3_io_ar_addr; // @[PHTS.scala 250:55]
  wire [2:0] PHTS_with_block_ram_3_io_ar_pht_addr; // @[PHTS.scala 250:55]
  wire [6:0] PHTS_with_block_ram_3_io_aw_addr; // @[PHTS.scala 250:55]
  wire [2:0] PHTS_with_block_ram_3_io_aw_pht_addr; // @[PHTS.scala 250:55]
  wire  PHTS_with_block_ram_3_io_write; // @[PHTS.scala 250:55]
  wire [7:0] PHTS_with_block_ram_3_io_in; // @[PHTS.scala 250:55]
  wire [7:0] PHTS_with_block_ram_3_io_pht_out; // @[PHTS.scala 250:55]
  wire [1:0] PHTS_with_block_ram_3_io_out; // @[PHTS.scala 250:55]
  reg [1:0] ar_bank_sel_reg; // @[PHTS.scala 261:34]
  wire [1:0] phts_banks_0_out = PHTS_with_block_ram_io_out; // @[PHTS.scala 250:{29,29}]
  wire [1:0] phts_banks_1_out = PHTS_with_block_ram_1_io_out; // @[PHTS.scala 250:{29,29}]
  wire [1:0] _GEN_1 = 2'h1 == ar_bank_sel_reg ? phts_banks_1_out : phts_banks_0_out; // @[PHTS.scala 263:{14,14}]
  wire [1:0] phts_banks_2_out = PHTS_with_block_ram_2_io_out; // @[PHTS.scala 250:{29,29}]
  wire [1:0] _GEN_2 = 2'h2 == ar_bank_sel_reg ? phts_banks_2_out : _GEN_1; // @[PHTS.scala 263:{14,14}]
  wire [1:0] phts_banks_3_out = PHTS_with_block_ram_3_io_out; // @[PHTS.scala 250:{29,29}]
  wire [7:0] phts_banks_0_pht_out = PHTS_with_block_ram_io_pht_out; // @[PHTS.scala 250:{29,29}]
  wire [7:0] phts_banks_1_pht_out = PHTS_with_block_ram_1_io_pht_out; // @[PHTS.scala 250:{29,29}]
  wire [7:0] _GEN_5 = 2'h1 == ar_bank_sel_reg ? phts_banks_1_pht_out : phts_banks_0_pht_out; // @[PHTS.scala 266:{16,16}]
  wire [7:0] phts_banks_2_pht_out = PHTS_with_block_ram_2_io_pht_out; // @[PHTS.scala 250:{29,29}]
  wire [7:0] _GEN_6 = 2'h2 == ar_bank_sel_reg ? phts_banks_2_pht_out : _GEN_5; // @[PHTS.scala 266:{16,16}]
  wire [7:0] phts_banks_3_pht_out = PHTS_with_block_ram_3_io_pht_out; // @[PHTS.scala 250:{29,29}]
  PHTS_with_block_ram PHTS_with_block_ram ( // @[PHTS.scala 250:55]
    .clock(PHTS_with_block_ram_clock),
    .reset(PHTS_with_block_ram_reset),
    .io_ar_addr(PHTS_with_block_ram_io_ar_addr),
    .io_ar_pht_addr(PHTS_with_block_ram_io_ar_pht_addr),
    .io_aw_addr(PHTS_with_block_ram_io_aw_addr),
    .io_aw_pht_addr(PHTS_with_block_ram_io_aw_pht_addr),
    .io_write(PHTS_with_block_ram_io_write),
    .io_in(PHTS_with_block_ram_io_in),
    .io_pht_out(PHTS_with_block_ram_io_pht_out),
    .io_out(PHTS_with_block_ram_io_out)
  );
  PHTS_with_block_ram PHTS_with_block_ram_1 ( // @[PHTS.scala 250:55]
    .clock(PHTS_with_block_ram_1_clock),
    .reset(PHTS_with_block_ram_1_reset),
    .io_ar_addr(PHTS_with_block_ram_1_io_ar_addr),
    .io_ar_pht_addr(PHTS_with_block_ram_1_io_ar_pht_addr),
    .io_aw_addr(PHTS_with_block_ram_1_io_aw_addr),
    .io_aw_pht_addr(PHTS_with_block_ram_1_io_aw_pht_addr),
    .io_write(PHTS_with_block_ram_1_io_write),
    .io_in(PHTS_with_block_ram_1_io_in),
    .io_pht_out(PHTS_with_block_ram_1_io_pht_out),
    .io_out(PHTS_with_block_ram_1_io_out)
  );
  PHTS_with_block_ram PHTS_with_block_ram_2 ( // @[PHTS.scala 250:55]
    .clock(PHTS_with_block_ram_2_clock),
    .reset(PHTS_with_block_ram_2_reset),
    .io_ar_addr(PHTS_with_block_ram_2_io_ar_addr),
    .io_ar_pht_addr(PHTS_with_block_ram_2_io_ar_pht_addr),
    .io_aw_addr(PHTS_with_block_ram_2_io_aw_addr),
    .io_aw_pht_addr(PHTS_with_block_ram_2_io_aw_pht_addr),
    .io_write(PHTS_with_block_ram_2_io_write),
    .io_in(PHTS_with_block_ram_2_io_in),
    .io_pht_out(PHTS_with_block_ram_2_io_pht_out),
    .io_out(PHTS_with_block_ram_2_io_out)
  );
  PHTS_with_block_ram PHTS_with_block_ram_3 ( // @[PHTS.scala 250:55]
    .clock(PHTS_with_block_ram_3_clock),
    .reset(PHTS_with_block_ram_3_reset),
    .io_ar_addr(PHTS_with_block_ram_3_io_ar_addr),
    .io_ar_pht_addr(PHTS_with_block_ram_3_io_ar_pht_addr),
    .io_aw_addr(PHTS_with_block_ram_3_io_aw_addr),
    .io_aw_pht_addr(PHTS_with_block_ram_3_io_aw_pht_addr),
    .io_write(PHTS_with_block_ram_3_io_write),
    .io_in(PHTS_with_block_ram_3_io_in),
    .io_pht_out(PHTS_with_block_ram_3_io_pht_out),
    .io_out(PHTS_with_block_ram_3_io_out)
  );
  assign io_out_L = 2'h3 == ar_bank_sel_reg ? phts_banks_3_out : _GEN_2; // @[PHTS.scala 263:{14,14}]
  assign io_pht_out = 2'h3 == ar_bank_sel_reg ? phts_banks_3_pht_out : _GEN_6; // @[PHTS.scala 266:{16,16}]
  assign PHTS_with_block_ram_clock = clock;
  assign PHTS_with_block_ram_reset = reset;
  assign PHTS_with_block_ram_io_ar_addr = io_ar_addr_L; // @[PHTS.scala 250:29 254:31]
  assign PHTS_with_block_ram_io_ar_pht_addr = io_ar_pht_addr; // @[PHTS.scala 250:29 257:35]
  assign PHTS_with_block_ram_io_aw_addr = io_aw_addr; // @[PHTS.scala 250:29 258:31]
  assign PHTS_with_block_ram_io_aw_pht_addr = io_aw_pht_addr; // @[PHTS.scala 250:29 259:35]
  assign PHTS_with_block_ram_io_write = io_aw_bank_sel == 2'h0 & io_write; // @[PHTS.scala 252:60]
  assign PHTS_with_block_ram_io_in = io_in; // @[PHTS.scala 250:29 253:26]
  assign PHTS_with_block_ram_1_clock = clock;
  assign PHTS_with_block_ram_1_reset = reset;
  assign PHTS_with_block_ram_1_io_ar_addr = io_ar_addr_L; // @[PHTS.scala 250:29 254:31]
  assign PHTS_with_block_ram_1_io_ar_pht_addr = io_ar_pht_addr; // @[PHTS.scala 250:29 257:35]
  assign PHTS_with_block_ram_1_io_aw_addr = io_aw_addr; // @[PHTS.scala 250:29 258:31]
  assign PHTS_with_block_ram_1_io_aw_pht_addr = io_aw_pht_addr; // @[PHTS.scala 250:29 259:35]
  assign PHTS_with_block_ram_1_io_write = io_aw_bank_sel == 2'h1 & io_write; // @[PHTS.scala 252:60]
  assign PHTS_with_block_ram_1_io_in = io_in; // @[PHTS.scala 250:29 253:26]
  assign PHTS_with_block_ram_2_clock = clock;
  assign PHTS_with_block_ram_2_reset = reset;
  assign PHTS_with_block_ram_2_io_ar_addr = io_ar_addr_L; // @[PHTS.scala 250:29 254:31]
  assign PHTS_with_block_ram_2_io_ar_pht_addr = io_ar_pht_addr; // @[PHTS.scala 250:29 257:35]
  assign PHTS_with_block_ram_2_io_aw_addr = io_aw_addr; // @[PHTS.scala 250:29 258:31]
  assign PHTS_with_block_ram_2_io_aw_pht_addr = io_aw_pht_addr; // @[PHTS.scala 250:29 259:35]
  assign PHTS_with_block_ram_2_io_write = io_aw_bank_sel == 2'h2 & io_write; // @[PHTS.scala 252:60]
  assign PHTS_with_block_ram_2_io_in = io_in; // @[PHTS.scala 250:29 253:26]
  assign PHTS_with_block_ram_3_clock = clock;
  assign PHTS_with_block_ram_3_reset = reset;
  assign PHTS_with_block_ram_3_io_ar_addr = io_ar_addr_L; // @[PHTS.scala 250:29 254:31]
  assign PHTS_with_block_ram_3_io_ar_pht_addr = io_ar_pht_addr; // @[PHTS.scala 250:29 257:35]
  assign PHTS_with_block_ram_3_io_aw_addr = io_aw_addr; // @[PHTS.scala 250:29 258:31]
  assign PHTS_with_block_ram_3_io_aw_pht_addr = io_aw_pht_addr; // @[PHTS.scala 250:29 259:35]
  assign PHTS_with_block_ram_3_io_write = io_aw_bank_sel == 2'h3 & io_write; // @[PHTS.scala 252:60]
  assign PHTS_with_block_ram_3_io_in = io_in; // @[PHTS.scala 250:29 253:26]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[PHTS.scala 261:34]
      ar_bank_sel_reg <= 2'h0; // @[PHTS.scala 261:34]
    end else begin
      ar_bank_sel_reg <= io_ar_bank_sel; // @[PHTS.scala 262:21]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ar_bank_sel_reg = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    ar_bank_sel_reg = 2'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BHT(
  input        clock,
  input        reset,
  input  [6:0] io_ar_addr,
  input  [6:0] io_aw_addr,
  input        io_write,
  input  [2:0] io_in,
  output [2:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] bht_0; // @[BHT.scala 20:22]
  reg [2:0] bht_1; // @[BHT.scala 20:22]
  reg [2:0] bht_2; // @[BHT.scala 20:22]
  reg [2:0] bht_3; // @[BHT.scala 20:22]
  reg [2:0] bht_4; // @[BHT.scala 20:22]
  reg [2:0] bht_5; // @[BHT.scala 20:22]
  reg [2:0] bht_6; // @[BHT.scala 20:22]
  reg [2:0] bht_7; // @[BHT.scala 20:22]
  reg [2:0] bht_8; // @[BHT.scala 20:22]
  reg [2:0] bht_9; // @[BHT.scala 20:22]
  reg [2:0] bht_10; // @[BHT.scala 20:22]
  reg [2:0] bht_11; // @[BHT.scala 20:22]
  reg [2:0] bht_12; // @[BHT.scala 20:22]
  reg [2:0] bht_13; // @[BHT.scala 20:22]
  reg [2:0] bht_14; // @[BHT.scala 20:22]
  reg [2:0] bht_15; // @[BHT.scala 20:22]
  reg [2:0] bht_16; // @[BHT.scala 20:22]
  reg [2:0] bht_17; // @[BHT.scala 20:22]
  reg [2:0] bht_18; // @[BHT.scala 20:22]
  reg [2:0] bht_19; // @[BHT.scala 20:22]
  reg [2:0] bht_20; // @[BHT.scala 20:22]
  reg [2:0] bht_21; // @[BHT.scala 20:22]
  reg [2:0] bht_22; // @[BHT.scala 20:22]
  reg [2:0] bht_23; // @[BHT.scala 20:22]
  reg [2:0] bht_24; // @[BHT.scala 20:22]
  reg [2:0] bht_25; // @[BHT.scala 20:22]
  reg [2:0] bht_26; // @[BHT.scala 20:22]
  reg [2:0] bht_27; // @[BHT.scala 20:22]
  reg [2:0] bht_28; // @[BHT.scala 20:22]
  reg [2:0] bht_29; // @[BHT.scala 20:22]
  reg [2:0] bht_30; // @[BHT.scala 20:22]
  reg [2:0] bht_31; // @[BHT.scala 20:22]
  reg [2:0] bht_32; // @[BHT.scala 20:22]
  reg [2:0] bht_33; // @[BHT.scala 20:22]
  reg [2:0] bht_34; // @[BHT.scala 20:22]
  reg [2:0] bht_35; // @[BHT.scala 20:22]
  reg [2:0] bht_36; // @[BHT.scala 20:22]
  reg [2:0] bht_37; // @[BHT.scala 20:22]
  reg [2:0] bht_38; // @[BHT.scala 20:22]
  reg [2:0] bht_39; // @[BHT.scala 20:22]
  reg [2:0] bht_40; // @[BHT.scala 20:22]
  reg [2:0] bht_41; // @[BHT.scala 20:22]
  reg [2:0] bht_42; // @[BHT.scala 20:22]
  reg [2:0] bht_43; // @[BHT.scala 20:22]
  reg [2:0] bht_44; // @[BHT.scala 20:22]
  reg [2:0] bht_45; // @[BHT.scala 20:22]
  reg [2:0] bht_46; // @[BHT.scala 20:22]
  reg [2:0] bht_47; // @[BHT.scala 20:22]
  reg [2:0] bht_48; // @[BHT.scala 20:22]
  reg [2:0] bht_49; // @[BHT.scala 20:22]
  reg [2:0] bht_50; // @[BHT.scala 20:22]
  reg [2:0] bht_51; // @[BHT.scala 20:22]
  reg [2:0] bht_52; // @[BHT.scala 20:22]
  reg [2:0] bht_53; // @[BHT.scala 20:22]
  reg [2:0] bht_54; // @[BHT.scala 20:22]
  reg [2:0] bht_55; // @[BHT.scala 20:22]
  reg [2:0] bht_56; // @[BHT.scala 20:22]
  reg [2:0] bht_57; // @[BHT.scala 20:22]
  reg [2:0] bht_58; // @[BHT.scala 20:22]
  reg [2:0] bht_59; // @[BHT.scala 20:22]
  reg [2:0] bht_60; // @[BHT.scala 20:22]
  reg [2:0] bht_61; // @[BHT.scala 20:22]
  reg [2:0] bht_62; // @[BHT.scala 20:22]
  reg [2:0] bht_63; // @[BHT.scala 20:22]
  reg [2:0] bht_64; // @[BHT.scala 20:22]
  reg [2:0] bht_65; // @[BHT.scala 20:22]
  reg [2:0] bht_66; // @[BHT.scala 20:22]
  reg [2:0] bht_67; // @[BHT.scala 20:22]
  reg [2:0] bht_68; // @[BHT.scala 20:22]
  reg [2:0] bht_69; // @[BHT.scala 20:22]
  reg [2:0] bht_70; // @[BHT.scala 20:22]
  reg [2:0] bht_71; // @[BHT.scala 20:22]
  reg [2:0] bht_72; // @[BHT.scala 20:22]
  reg [2:0] bht_73; // @[BHT.scala 20:22]
  reg [2:0] bht_74; // @[BHT.scala 20:22]
  reg [2:0] bht_75; // @[BHT.scala 20:22]
  reg [2:0] bht_76; // @[BHT.scala 20:22]
  reg [2:0] bht_77; // @[BHT.scala 20:22]
  reg [2:0] bht_78; // @[BHT.scala 20:22]
  reg [2:0] bht_79; // @[BHT.scala 20:22]
  reg [2:0] bht_80; // @[BHT.scala 20:22]
  reg [2:0] bht_81; // @[BHT.scala 20:22]
  reg [2:0] bht_82; // @[BHT.scala 20:22]
  reg [2:0] bht_83; // @[BHT.scala 20:22]
  reg [2:0] bht_84; // @[BHT.scala 20:22]
  reg [2:0] bht_85; // @[BHT.scala 20:22]
  reg [2:0] bht_86; // @[BHT.scala 20:22]
  reg [2:0] bht_87; // @[BHT.scala 20:22]
  reg [2:0] bht_88; // @[BHT.scala 20:22]
  reg [2:0] bht_89; // @[BHT.scala 20:22]
  reg [2:0] bht_90; // @[BHT.scala 20:22]
  reg [2:0] bht_91; // @[BHT.scala 20:22]
  reg [2:0] bht_92; // @[BHT.scala 20:22]
  reg [2:0] bht_93; // @[BHT.scala 20:22]
  reg [2:0] bht_94; // @[BHT.scala 20:22]
  reg [2:0] bht_95; // @[BHT.scala 20:22]
  reg [2:0] bht_96; // @[BHT.scala 20:22]
  reg [2:0] bht_97; // @[BHT.scala 20:22]
  reg [2:0] bht_98; // @[BHT.scala 20:22]
  reg [2:0] bht_99; // @[BHT.scala 20:22]
  reg [2:0] bht_100; // @[BHT.scala 20:22]
  reg [2:0] bht_101; // @[BHT.scala 20:22]
  reg [2:0] bht_102; // @[BHT.scala 20:22]
  reg [2:0] bht_103; // @[BHT.scala 20:22]
  reg [2:0] bht_104; // @[BHT.scala 20:22]
  reg [2:0] bht_105; // @[BHT.scala 20:22]
  reg [2:0] bht_106; // @[BHT.scala 20:22]
  reg [2:0] bht_107; // @[BHT.scala 20:22]
  reg [2:0] bht_108; // @[BHT.scala 20:22]
  reg [2:0] bht_109; // @[BHT.scala 20:22]
  reg [2:0] bht_110; // @[BHT.scala 20:22]
  reg [2:0] bht_111; // @[BHT.scala 20:22]
  reg [2:0] bht_112; // @[BHT.scala 20:22]
  reg [2:0] bht_113; // @[BHT.scala 20:22]
  reg [2:0] bht_114; // @[BHT.scala 20:22]
  reg [2:0] bht_115; // @[BHT.scala 20:22]
  reg [2:0] bht_116; // @[BHT.scala 20:22]
  reg [2:0] bht_117; // @[BHT.scala 20:22]
  reg [2:0] bht_118; // @[BHT.scala 20:22]
  reg [2:0] bht_119; // @[BHT.scala 20:22]
  reg [2:0] bht_120; // @[BHT.scala 20:22]
  reg [2:0] bht_121; // @[BHT.scala 20:22]
  reg [2:0] bht_122; // @[BHT.scala 20:22]
  reg [2:0] bht_123; // @[BHT.scala 20:22]
  reg [2:0] bht_124; // @[BHT.scala 20:22]
  reg [2:0] bht_125; // @[BHT.scala 20:22]
  reg [2:0] bht_126; // @[BHT.scala 20:22]
  reg [2:0] bht_127; // @[BHT.scala 20:22]
  wire [2:0] _GEN_1 = 7'h1 == io_ar_addr ? bht_1 : bht_0; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_2 = 7'h2 == io_ar_addr ? bht_2 : _GEN_1; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_3 = 7'h3 == io_ar_addr ? bht_3 : _GEN_2; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_4 = 7'h4 == io_ar_addr ? bht_4 : _GEN_3; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_5 = 7'h5 == io_ar_addr ? bht_5 : _GEN_4; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_6 = 7'h6 == io_ar_addr ? bht_6 : _GEN_5; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_7 = 7'h7 == io_ar_addr ? bht_7 : _GEN_6; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_8 = 7'h8 == io_ar_addr ? bht_8 : _GEN_7; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_9 = 7'h9 == io_ar_addr ? bht_9 : _GEN_8; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_10 = 7'ha == io_ar_addr ? bht_10 : _GEN_9; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_11 = 7'hb == io_ar_addr ? bht_11 : _GEN_10; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_12 = 7'hc == io_ar_addr ? bht_12 : _GEN_11; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_13 = 7'hd == io_ar_addr ? bht_13 : _GEN_12; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_14 = 7'he == io_ar_addr ? bht_14 : _GEN_13; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_15 = 7'hf == io_ar_addr ? bht_15 : _GEN_14; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_16 = 7'h10 == io_ar_addr ? bht_16 : _GEN_15; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_17 = 7'h11 == io_ar_addr ? bht_17 : _GEN_16; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_18 = 7'h12 == io_ar_addr ? bht_18 : _GEN_17; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_19 = 7'h13 == io_ar_addr ? bht_19 : _GEN_18; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_20 = 7'h14 == io_ar_addr ? bht_20 : _GEN_19; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_21 = 7'h15 == io_ar_addr ? bht_21 : _GEN_20; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_22 = 7'h16 == io_ar_addr ? bht_22 : _GEN_21; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_23 = 7'h17 == io_ar_addr ? bht_23 : _GEN_22; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_24 = 7'h18 == io_ar_addr ? bht_24 : _GEN_23; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_25 = 7'h19 == io_ar_addr ? bht_25 : _GEN_24; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_26 = 7'h1a == io_ar_addr ? bht_26 : _GEN_25; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_27 = 7'h1b == io_ar_addr ? bht_27 : _GEN_26; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_28 = 7'h1c == io_ar_addr ? bht_28 : _GEN_27; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_29 = 7'h1d == io_ar_addr ? bht_29 : _GEN_28; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_30 = 7'h1e == io_ar_addr ? bht_30 : _GEN_29; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_31 = 7'h1f == io_ar_addr ? bht_31 : _GEN_30; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_32 = 7'h20 == io_ar_addr ? bht_32 : _GEN_31; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_33 = 7'h21 == io_ar_addr ? bht_33 : _GEN_32; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_34 = 7'h22 == io_ar_addr ? bht_34 : _GEN_33; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_35 = 7'h23 == io_ar_addr ? bht_35 : _GEN_34; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_36 = 7'h24 == io_ar_addr ? bht_36 : _GEN_35; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_37 = 7'h25 == io_ar_addr ? bht_37 : _GEN_36; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_38 = 7'h26 == io_ar_addr ? bht_38 : _GEN_37; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_39 = 7'h27 == io_ar_addr ? bht_39 : _GEN_38; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_40 = 7'h28 == io_ar_addr ? bht_40 : _GEN_39; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_41 = 7'h29 == io_ar_addr ? bht_41 : _GEN_40; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_42 = 7'h2a == io_ar_addr ? bht_42 : _GEN_41; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_43 = 7'h2b == io_ar_addr ? bht_43 : _GEN_42; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_44 = 7'h2c == io_ar_addr ? bht_44 : _GEN_43; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_45 = 7'h2d == io_ar_addr ? bht_45 : _GEN_44; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_46 = 7'h2e == io_ar_addr ? bht_46 : _GEN_45; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_47 = 7'h2f == io_ar_addr ? bht_47 : _GEN_46; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_48 = 7'h30 == io_ar_addr ? bht_48 : _GEN_47; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_49 = 7'h31 == io_ar_addr ? bht_49 : _GEN_48; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_50 = 7'h32 == io_ar_addr ? bht_50 : _GEN_49; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_51 = 7'h33 == io_ar_addr ? bht_51 : _GEN_50; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_52 = 7'h34 == io_ar_addr ? bht_52 : _GEN_51; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_53 = 7'h35 == io_ar_addr ? bht_53 : _GEN_52; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_54 = 7'h36 == io_ar_addr ? bht_54 : _GEN_53; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_55 = 7'h37 == io_ar_addr ? bht_55 : _GEN_54; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_56 = 7'h38 == io_ar_addr ? bht_56 : _GEN_55; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_57 = 7'h39 == io_ar_addr ? bht_57 : _GEN_56; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_58 = 7'h3a == io_ar_addr ? bht_58 : _GEN_57; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_59 = 7'h3b == io_ar_addr ? bht_59 : _GEN_58; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_60 = 7'h3c == io_ar_addr ? bht_60 : _GEN_59; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_61 = 7'h3d == io_ar_addr ? bht_61 : _GEN_60; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_62 = 7'h3e == io_ar_addr ? bht_62 : _GEN_61; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_63 = 7'h3f == io_ar_addr ? bht_63 : _GEN_62; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_64 = 7'h40 == io_ar_addr ? bht_64 : _GEN_63; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_65 = 7'h41 == io_ar_addr ? bht_65 : _GEN_64; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_66 = 7'h42 == io_ar_addr ? bht_66 : _GEN_65; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_67 = 7'h43 == io_ar_addr ? bht_67 : _GEN_66; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_68 = 7'h44 == io_ar_addr ? bht_68 : _GEN_67; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_69 = 7'h45 == io_ar_addr ? bht_69 : _GEN_68; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_70 = 7'h46 == io_ar_addr ? bht_70 : _GEN_69; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_71 = 7'h47 == io_ar_addr ? bht_71 : _GEN_70; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_72 = 7'h48 == io_ar_addr ? bht_72 : _GEN_71; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_73 = 7'h49 == io_ar_addr ? bht_73 : _GEN_72; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_74 = 7'h4a == io_ar_addr ? bht_74 : _GEN_73; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_75 = 7'h4b == io_ar_addr ? bht_75 : _GEN_74; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_76 = 7'h4c == io_ar_addr ? bht_76 : _GEN_75; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_77 = 7'h4d == io_ar_addr ? bht_77 : _GEN_76; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_78 = 7'h4e == io_ar_addr ? bht_78 : _GEN_77; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_79 = 7'h4f == io_ar_addr ? bht_79 : _GEN_78; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_80 = 7'h50 == io_ar_addr ? bht_80 : _GEN_79; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_81 = 7'h51 == io_ar_addr ? bht_81 : _GEN_80; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_82 = 7'h52 == io_ar_addr ? bht_82 : _GEN_81; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_83 = 7'h53 == io_ar_addr ? bht_83 : _GEN_82; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_84 = 7'h54 == io_ar_addr ? bht_84 : _GEN_83; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_85 = 7'h55 == io_ar_addr ? bht_85 : _GEN_84; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_86 = 7'h56 == io_ar_addr ? bht_86 : _GEN_85; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_87 = 7'h57 == io_ar_addr ? bht_87 : _GEN_86; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_88 = 7'h58 == io_ar_addr ? bht_88 : _GEN_87; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_89 = 7'h59 == io_ar_addr ? bht_89 : _GEN_88; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_90 = 7'h5a == io_ar_addr ? bht_90 : _GEN_89; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_91 = 7'h5b == io_ar_addr ? bht_91 : _GEN_90; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_92 = 7'h5c == io_ar_addr ? bht_92 : _GEN_91; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_93 = 7'h5d == io_ar_addr ? bht_93 : _GEN_92; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_94 = 7'h5e == io_ar_addr ? bht_94 : _GEN_93; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_95 = 7'h5f == io_ar_addr ? bht_95 : _GEN_94; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_96 = 7'h60 == io_ar_addr ? bht_96 : _GEN_95; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_97 = 7'h61 == io_ar_addr ? bht_97 : _GEN_96; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_98 = 7'h62 == io_ar_addr ? bht_98 : _GEN_97; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_99 = 7'h63 == io_ar_addr ? bht_99 : _GEN_98; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_100 = 7'h64 == io_ar_addr ? bht_100 : _GEN_99; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_101 = 7'h65 == io_ar_addr ? bht_101 : _GEN_100; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_102 = 7'h66 == io_ar_addr ? bht_102 : _GEN_101; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_103 = 7'h67 == io_ar_addr ? bht_103 : _GEN_102; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_104 = 7'h68 == io_ar_addr ? bht_104 : _GEN_103; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_105 = 7'h69 == io_ar_addr ? bht_105 : _GEN_104; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_106 = 7'h6a == io_ar_addr ? bht_106 : _GEN_105; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_107 = 7'h6b == io_ar_addr ? bht_107 : _GEN_106; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_108 = 7'h6c == io_ar_addr ? bht_108 : _GEN_107; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_109 = 7'h6d == io_ar_addr ? bht_109 : _GEN_108; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_110 = 7'h6e == io_ar_addr ? bht_110 : _GEN_109; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_111 = 7'h6f == io_ar_addr ? bht_111 : _GEN_110; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_112 = 7'h70 == io_ar_addr ? bht_112 : _GEN_111; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_113 = 7'h71 == io_ar_addr ? bht_113 : _GEN_112; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_114 = 7'h72 == io_ar_addr ? bht_114 : _GEN_113; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_115 = 7'h73 == io_ar_addr ? bht_115 : _GEN_114; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_116 = 7'h74 == io_ar_addr ? bht_116 : _GEN_115; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_117 = 7'h75 == io_ar_addr ? bht_117 : _GEN_116; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_118 = 7'h76 == io_ar_addr ? bht_118 : _GEN_117; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_119 = 7'h77 == io_ar_addr ? bht_119 : _GEN_118; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_120 = 7'h78 == io_ar_addr ? bht_120 : _GEN_119; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_121 = 7'h79 == io_ar_addr ? bht_121 : _GEN_120; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_122 = 7'h7a == io_ar_addr ? bht_122 : _GEN_121; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_123 = 7'h7b == io_ar_addr ? bht_123 : _GEN_122; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_124 = 7'h7c == io_ar_addr ? bht_124 : _GEN_123; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_125 = 7'h7d == io_ar_addr ? bht_125 : _GEN_124; // @[BHT.scala 21:{12,12}]
  wire [2:0] _GEN_126 = 7'h7e == io_ar_addr ? bht_126 : _GEN_125; // @[BHT.scala 21:{12,12}]
  assign io_out = 7'h7f == io_ar_addr ? bht_127 : _GEN_126; // @[BHT.scala 21:{12,12}]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_0 <= 3'h0;
    end else if (io_write & 7'h0 == io_aw_addr) begin
      bht_0 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_1 <= 3'h0;
    end else if (io_write & 7'h1 == io_aw_addr) begin
      bht_1 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_2 <= 3'h0;
    end else if (io_write & 7'h2 == io_aw_addr) begin
      bht_2 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_3 <= 3'h0;
    end else if (io_write & 7'h3 == io_aw_addr) begin
      bht_3 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_4 <= 3'h0;
    end else if (io_write & 7'h4 == io_aw_addr) begin
      bht_4 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_5 <= 3'h0;
    end else if (io_write & 7'h5 == io_aw_addr) begin
      bht_5 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_6 <= 3'h0;
    end else if (io_write & 7'h6 == io_aw_addr) begin
      bht_6 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_7 <= 3'h0;
    end else if (io_write & 7'h7 == io_aw_addr) begin
      bht_7 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_8 <= 3'h0;
    end else if (io_write & 7'h8 == io_aw_addr) begin
      bht_8 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_9 <= 3'h0;
    end else if (io_write & 7'h9 == io_aw_addr) begin
      bht_9 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_10 <= 3'h0;
    end else if (io_write & 7'ha == io_aw_addr) begin
      bht_10 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_11 <= 3'h0;
    end else if (io_write & 7'hb == io_aw_addr) begin
      bht_11 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_12 <= 3'h0;
    end else if (io_write & 7'hc == io_aw_addr) begin
      bht_12 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_13 <= 3'h0;
    end else if (io_write & 7'hd == io_aw_addr) begin
      bht_13 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_14 <= 3'h0;
    end else if (io_write & 7'he == io_aw_addr) begin
      bht_14 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_15 <= 3'h0;
    end else if (io_write & 7'hf == io_aw_addr) begin
      bht_15 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_16 <= 3'h0;
    end else if (io_write & 7'h10 == io_aw_addr) begin
      bht_16 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_17 <= 3'h0;
    end else if (io_write & 7'h11 == io_aw_addr) begin
      bht_17 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_18 <= 3'h0;
    end else if (io_write & 7'h12 == io_aw_addr) begin
      bht_18 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_19 <= 3'h0;
    end else if (io_write & 7'h13 == io_aw_addr) begin
      bht_19 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_20 <= 3'h0;
    end else if (io_write & 7'h14 == io_aw_addr) begin
      bht_20 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_21 <= 3'h0;
    end else if (io_write & 7'h15 == io_aw_addr) begin
      bht_21 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_22 <= 3'h0;
    end else if (io_write & 7'h16 == io_aw_addr) begin
      bht_22 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_23 <= 3'h0;
    end else if (io_write & 7'h17 == io_aw_addr) begin
      bht_23 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_24 <= 3'h0;
    end else if (io_write & 7'h18 == io_aw_addr) begin
      bht_24 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_25 <= 3'h0;
    end else if (io_write & 7'h19 == io_aw_addr) begin
      bht_25 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_26 <= 3'h0;
    end else if (io_write & 7'h1a == io_aw_addr) begin
      bht_26 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_27 <= 3'h0;
    end else if (io_write & 7'h1b == io_aw_addr) begin
      bht_27 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_28 <= 3'h0;
    end else if (io_write & 7'h1c == io_aw_addr) begin
      bht_28 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_29 <= 3'h0;
    end else if (io_write & 7'h1d == io_aw_addr) begin
      bht_29 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_30 <= 3'h0;
    end else if (io_write & 7'h1e == io_aw_addr) begin
      bht_30 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_31 <= 3'h0;
    end else if (io_write & 7'h1f == io_aw_addr) begin
      bht_31 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_32 <= 3'h0;
    end else if (io_write & 7'h20 == io_aw_addr) begin
      bht_32 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_33 <= 3'h0;
    end else if (io_write & 7'h21 == io_aw_addr) begin
      bht_33 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_34 <= 3'h0;
    end else if (io_write & 7'h22 == io_aw_addr) begin
      bht_34 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_35 <= 3'h0;
    end else if (io_write & 7'h23 == io_aw_addr) begin
      bht_35 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_36 <= 3'h0;
    end else if (io_write & 7'h24 == io_aw_addr) begin
      bht_36 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_37 <= 3'h0;
    end else if (io_write & 7'h25 == io_aw_addr) begin
      bht_37 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_38 <= 3'h0;
    end else if (io_write & 7'h26 == io_aw_addr) begin
      bht_38 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_39 <= 3'h0;
    end else if (io_write & 7'h27 == io_aw_addr) begin
      bht_39 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_40 <= 3'h0;
    end else if (io_write & 7'h28 == io_aw_addr) begin
      bht_40 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_41 <= 3'h0;
    end else if (io_write & 7'h29 == io_aw_addr) begin
      bht_41 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_42 <= 3'h0;
    end else if (io_write & 7'h2a == io_aw_addr) begin
      bht_42 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_43 <= 3'h0;
    end else if (io_write & 7'h2b == io_aw_addr) begin
      bht_43 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_44 <= 3'h0;
    end else if (io_write & 7'h2c == io_aw_addr) begin
      bht_44 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_45 <= 3'h0;
    end else if (io_write & 7'h2d == io_aw_addr) begin
      bht_45 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_46 <= 3'h0;
    end else if (io_write & 7'h2e == io_aw_addr) begin
      bht_46 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_47 <= 3'h0;
    end else if (io_write & 7'h2f == io_aw_addr) begin
      bht_47 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_48 <= 3'h0;
    end else if (io_write & 7'h30 == io_aw_addr) begin
      bht_48 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_49 <= 3'h0;
    end else if (io_write & 7'h31 == io_aw_addr) begin
      bht_49 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_50 <= 3'h0;
    end else if (io_write & 7'h32 == io_aw_addr) begin
      bht_50 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_51 <= 3'h0;
    end else if (io_write & 7'h33 == io_aw_addr) begin
      bht_51 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_52 <= 3'h0;
    end else if (io_write & 7'h34 == io_aw_addr) begin
      bht_52 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_53 <= 3'h0;
    end else if (io_write & 7'h35 == io_aw_addr) begin
      bht_53 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_54 <= 3'h0;
    end else if (io_write & 7'h36 == io_aw_addr) begin
      bht_54 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_55 <= 3'h0;
    end else if (io_write & 7'h37 == io_aw_addr) begin
      bht_55 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_56 <= 3'h0;
    end else if (io_write & 7'h38 == io_aw_addr) begin
      bht_56 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_57 <= 3'h0;
    end else if (io_write & 7'h39 == io_aw_addr) begin
      bht_57 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_58 <= 3'h0;
    end else if (io_write & 7'h3a == io_aw_addr) begin
      bht_58 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_59 <= 3'h0;
    end else if (io_write & 7'h3b == io_aw_addr) begin
      bht_59 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_60 <= 3'h0;
    end else if (io_write & 7'h3c == io_aw_addr) begin
      bht_60 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_61 <= 3'h0;
    end else if (io_write & 7'h3d == io_aw_addr) begin
      bht_61 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_62 <= 3'h0;
    end else if (io_write & 7'h3e == io_aw_addr) begin
      bht_62 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_63 <= 3'h0;
    end else if (io_write & 7'h3f == io_aw_addr) begin
      bht_63 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_64 <= 3'h0;
    end else if (io_write & 7'h40 == io_aw_addr) begin
      bht_64 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_65 <= 3'h0;
    end else if (io_write & 7'h41 == io_aw_addr) begin
      bht_65 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_66 <= 3'h0;
    end else if (io_write & 7'h42 == io_aw_addr) begin
      bht_66 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_67 <= 3'h0;
    end else if (io_write & 7'h43 == io_aw_addr) begin
      bht_67 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_68 <= 3'h0;
    end else if (io_write & 7'h44 == io_aw_addr) begin
      bht_68 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_69 <= 3'h0;
    end else if (io_write & 7'h45 == io_aw_addr) begin
      bht_69 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_70 <= 3'h0;
    end else if (io_write & 7'h46 == io_aw_addr) begin
      bht_70 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_71 <= 3'h0;
    end else if (io_write & 7'h47 == io_aw_addr) begin
      bht_71 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_72 <= 3'h0;
    end else if (io_write & 7'h48 == io_aw_addr) begin
      bht_72 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_73 <= 3'h0;
    end else if (io_write & 7'h49 == io_aw_addr) begin
      bht_73 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_74 <= 3'h0;
    end else if (io_write & 7'h4a == io_aw_addr) begin
      bht_74 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_75 <= 3'h0;
    end else if (io_write & 7'h4b == io_aw_addr) begin
      bht_75 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_76 <= 3'h0;
    end else if (io_write & 7'h4c == io_aw_addr) begin
      bht_76 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_77 <= 3'h0;
    end else if (io_write & 7'h4d == io_aw_addr) begin
      bht_77 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_78 <= 3'h0;
    end else if (io_write & 7'h4e == io_aw_addr) begin
      bht_78 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_79 <= 3'h0;
    end else if (io_write & 7'h4f == io_aw_addr) begin
      bht_79 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_80 <= 3'h0;
    end else if (io_write & 7'h50 == io_aw_addr) begin
      bht_80 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_81 <= 3'h0;
    end else if (io_write & 7'h51 == io_aw_addr) begin
      bht_81 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_82 <= 3'h0;
    end else if (io_write & 7'h52 == io_aw_addr) begin
      bht_82 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_83 <= 3'h0;
    end else if (io_write & 7'h53 == io_aw_addr) begin
      bht_83 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_84 <= 3'h0;
    end else if (io_write & 7'h54 == io_aw_addr) begin
      bht_84 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_85 <= 3'h0;
    end else if (io_write & 7'h55 == io_aw_addr) begin
      bht_85 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_86 <= 3'h0;
    end else if (io_write & 7'h56 == io_aw_addr) begin
      bht_86 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_87 <= 3'h0;
    end else if (io_write & 7'h57 == io_aw_addr) begin
      bht_87 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_88 <= 3'h0;
    end else if (io_write & 7'h58 == io_aw_addr) begin
      bht_88 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_89 <= 3'h0;
    end else if (io_write & 7'h59 == io_aw_addr) begin
      bht_89 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_90 <= 3'h0;
    end else if (io_write & 7'h5a == io_aw_addr) begin
      bht_90 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_91 <= 3'h0;
    end else if (io_write & 7'h5b == io_aw_addr) begin
      bht_91 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_92 <= 3'h0;
    end else if (io_write & 7'h5c == io_aw_addr) begin
      bht_92 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_93 <= 3'h0;
    end else if (io_write & 7'h5d == io_aw_addr) begin
      bht_93 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_94 <= 3'h0;
    end else if (io_write & 7'h5e == io_aw_addr) begin
      bht_94 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_95 <= 3'h0;
    end else if (io_write & 7'h5f == io_aw_addr) begin
      bht_95 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_96 <= 3'h0;
    end else if (io_write & 7'h60 == io_aw_addr) begin
      bht_96 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_97 <= 3'h0;
    end else if (io_write & 7'h61 == io_aw_addr) begin
      bht_97 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_98 <= 3'h0;
    end else if (io_write & 7'h62 == io_aw_addr) begin
      bht_98 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_99 <= 3'h0;
    end else if (io_write & 7'h63 == io_aw_addr) begin
      bht_99 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_100 <= 3'h0;
    end else if (io_write & 7'h64 == io_aw_addr) begin
      bht_100 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_101 <= 3'h0;
    end else if (io_write & 7'h65 == io_aw_addr) begin
      bht_101 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_102 <= 3'h0;
    end else if (io_write & 7'h66 == io_aw_addr) begin
      bht_102 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_103 <= 3'h0;
    end else if (io_write & 7'h67 == io_aw_addr) begin
      bht_103 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_104 <= 3'h0;
    end else if (io_write & 7'h68 == io_aw_addr) begin
      bht_104 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_105 <= 3'h0;
    end else if (io_write & 7'h69 == io_aw_addr) begin
      bht_105 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_106 <= 3'h0;
    end else if (io_write & 7'h6a == io_aw_addr) begin
      bht_106 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_107 <= 3'h0;
    end else if (io_write & 7'h6b == io_aw_addr) begin
      bht_107 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_108 <= 3'h0;
    end else if (io_write & 7'h6c == io_aw_addr) begin
      bht_108 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_109 <= 3'h0;
    end else if (io_write & 7'h6d == io_aw_addr) begin
      bht_109 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_110 <= 3'h0;
    end else if (io_write & 7'h6e == io_aw_addr) begin
      bht_110 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_111 <= 3'h0;
    end else if (io_write & 7'h6f == io_aw_addr) begin
      bht_111 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_112 <= 3'h0;
    end else if (io_write & 7'h70 == io_aw_addr) begin
      bht_112 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_113 <= 3'h0;
    end else if (io_write & 7'h71 == io_aw_addr) begin
      bht_113 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_114 <= 3'h0;
    end else if (io_write & 7'h72 == io_aw_addr) begin
      bht_114 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_115 <= 3'h0;
    end else if (io_write & 7'h73 == io_aw_addr) begin
      bht_115 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_116 <= 3'h0;
    end else if (io_write & 7'h74 == io_aw_addr) begin
      bht_116 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_117 <= 3'h0;
    end else if (io_write & 7'h75 == io_aw_addr) begin
      bht_117 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_118 <= 3'h0;
    end else if (io_write & 7'h76 == io_aw_addr) begin
      bht_118 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_119 <= 3'h0;
    end else if (io_write & 7'h77 == io_aw_addr) begin
      bht_119 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_120 <= 3'h0;
    end else if (io_write & 7'h78 == io_aw_addr) begin
      bht_120 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_121 <= 3'h0;
    end else if (io_write & 7'h79 == io_aw_addr) begin
      bht_121 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_122 <= 3'h0;
    end else if (io_write & 7'h7a == io_aw_addr) begin
      bht_122 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_123 <= 3'h0;
    end else if (io_write & 7'h7b == io_aw_addr) begin
      bht_123 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_124 <= 3'h0;
    end else if (io_write & 7'h7c == io_aw_addr) begin
      bht_124 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_125 <= 3'h0;
    end else if (io_write & 7'h7d == io_aw_addr) begin
      bht_125 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_126 <= 3'h0;
    end else if (io_write & 7'h7e == io_aw_addr) begin
      bht_126 <= io_in;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BHT.scala 23:22]
      bht_127 <= 3'h0;
    end else if (io_write & 7'h7f == io_aw_addr) begin
      bht_127 <= io_in;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  bht_0 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  bht_1 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  bht_2 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  bht_3 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  bht_4 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  bht_5 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  bht_6 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  bht_7 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  bht_8 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  bht_9 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  bht_10 = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  bht_11 = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  bht_12 = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  bht_13 = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  bht_14 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  bht_15 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  bht_16 = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  bht_17 = _RAND_17[2:0];
  _RAND_18 = {1{`RANDOM}};
  bht_18 = _RAND_18[2:0];
  _RAND_19 = {1{`RANDOM}};
  bht_19 = _RAND_19[2:0];
  _RAND_20 = {1{`RANDOM}};
  bht_20 = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  bht_21 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  bht_22 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  bht_23 = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  bht_24 = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  bht_25 = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  bht_26 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  bht_27 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  bht_28 = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  bht_29 = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  bht_30 = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  bht_31 = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  bht_32 = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  bht_33 = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  bht_34 = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  bht_35 = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  bht_36 = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  bht_37 = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  bht_38 = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  bht_39 = _RAND_39[2:0];
  _RAND_40 = {1{`RANDOM}};
  bht_40 = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  bht_41 = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  bht_42 = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  bht_43 = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  bht_44 = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  bht_45 = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  bht_46 = _RAND_46[2:0];
  _RAND_47 = {1{`RANDOM}};
  bht_47 = _RAND_47[2:0];
  _RAND_48 = {1{`RANDOM}};
  bht_48 = _RAND_48[2:0];
  _RAND_49 = {1{`RANDOM}};
  bht_49 = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  bht_50 = _RAND_50[2:0];
  _RAND_51 = {1{`RANDOM}};
  bht_51 = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  bht_52 = _RAND_52[2:0];
  _RAND_53 = {1{`RANDOM}};
  bht_53 = _RAND_53[2:0];
  _RAND_54 = {1{`RANDOM}};
  bht_54 = _RAND_54[2:0];
  _RAND_55 = {1{`RANDOM}};
  bht_55 = _RAND_55[2:0];
  _RAND_56 = {1{`RANDOM}};
  bht_56 = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  bht_57 = _RAND_57[2:0];
  _RAND_58 = {1{`RANDOM}};
  bht_58 = _RAND_58[2:0];
  _RAND_59 = {1{`RANDOM}};
  bht_59 = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  bht_60 = _RAND_60[2:0];
  _RAND_61 = {1{`RANDOM}};
  bht_61 = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  bht_62 = _RAND_62[2:0];
  _RAND_63 = {1{`RANDOM}};
  bht_63 = _RAND_63[2:0];
  _RAND_64 = {1{`RANDOM}};
  bht_64 = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  bht_65 = _RAND_65[2:0];
  _RAND_66 = {1{`RANDOM}};
  bht_66 = _RAND_66[2:0];
  _RAND_67 = {1{`RANDOM}};
  bht_67 = _RAND_67[2:0];
  _RAND_68 = {1{`RANDOM}};
  bht_68 = _RAND_68[2:0];
  _RAND_69 = {1{`RANDOM}};
  bht_69 = _RAND_69[2:0];
  _RAND_70 = {1{`RANDOM}};
  bht_70 = _RAND_70[2:0];
  _RAND_71 = {1{`RANDOM}};
  bht_71 = _RAND_71[2:0];
  _RAND_72 = {1{`RANDOM}};
  bht_72 = _RAND_72[2:0];
  _RAND_73 = {1{`RANDOM}};
  bht_73 = _RAND_73[2:0];
  _RAND_74 = {1{`RANDOM}};
  bht_74 = _RAND_74[2:0];
  _RAND_75 = {1{`RANDOM}};
  bht_75 = _RAND_75[2:0];
  _RAND_76 = {1{`RANDOM}};
  bht_76 = _RAND_76[2:0];
  _RAND_77 = {1{`RANDOM}};
  bht_77 = _RAND_77[2:0];
  _RAND_78 = {1{`RANDOM}};
  bht_78 = _RAND_78[2:0];
  _RAND_79 = {1{`RANDOM}};
  bht_79 = _RAND_79[2:0];
  _RAND_80 = {1{`RANDOM}};
  bht_80 = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  bht_81 = _RAND_81[2:0];
  _RAND_82 = {1{`RANDOM}};
  bht_82 = _RAND_82[2:0];
  _RAND_83 = {1{`RANDOM}};
  bht_83 = _RAND_83[2:0];
  _RAND_84 = {1{`RANDOM}};
  bht_84 = _RAND_84[2:0];
  _RAND_85 = {1{`RANDOM}};
  bht_85 = _RAND_85[2:0];
  _RAND_86 = {1{`RANDOM}};
  bht_86 = _RAND_86[2:0];
  _RAND_87 = {1{`RANDOM}};
  bht_87 = _RAND_87[2:0];
  _RAND_88 = {1{`RANDOM}};
  bht_88 = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  bht_89 = _RAND_89[2:0];
  _RAND_90 = {1{`RANDOM}};
  bht_90 = _RAND_90[2:0];
  _RAND_91 = {1{`RANDOM}};
  bht_91 = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  bht_92 = _RAND_92[2:0];
  _RAND_93 = {1{`RANDOM}};
  bht_93 = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  bht_94 = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  bht_95 = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  bht_96 = _RAND_96[2:0];
  _RAND_97 = {1{`RANDOM}};
  bht_97 = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  bht_98 = _RAND_98[2:0];
  _RAND_99 = {1{`RANDOM}};
  bht_99 = _RAND_99[2:0];
  _RAND_100 = {1{`RANDOM}};
  bht_100 = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  bht_101 = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  bht_102 = _RAND_102[2:0];
  _RAND_103 = {1{`RANDOM}};
  bht_103 = _RAND_103[2:0];
  _RAND_104 = {1{`RANDOM}};
  bht_104 = _RAND_104[2:0];
  _RAND_105 = {1{`RANDOM}};
  bht_105 = _RAND_105[2:0];
  _RAND_106 = {1{`RANDOM}};
  bht_106 = _RAND_106[2:0];
  _RAND_107 = {1{`RANDOM}};
  bht_107 = _RAND_107[2:0];
  _RAND_108 = {1{`RANDOM}};
  bht_108 = _RAND_108[2:0];
  _RAND_109 = {1{`RANDOM}};
  bht_109 = _RAND_109[2:0];
  _RAND_110 = {1{`RANDOM}};
  bht_110 = _RAND_110[2:0];
  _RAND_111 = {1{`RANDOM}};
  bht_111 = _RAND_111[2:0];
  _RAND_112 = {1{`RANDOM}};
  bht_112 = _RAND_112[2:0];
  _RAND_113 = {1{`RANDOM}};
  bht_113 = _RAND_113[2:0];
  _RAND_114 = {1{`RANDOM}};
  bht_114 = _RAND_114[2:0];
  _RAND_115 = {1{`RANDOM}};
  bht_115 = _RAND_115[2:0];
  _RAND_116 = {1{`RANDOM}};
  bht_116 = _RAND_116[2:0];
  _RAND_117 = {1{`RANDOM}};
  bht_117 = _RAND_117[2:0];
  _RAND_118 = {1{`RANDOM}};
  bht_118 = _RAND_118[2:0];
  _RAND_119 = {1{`RANDOM}};
  bht_119 = _RAND_119[2:0];
  _RAND_120 = {1{`RANDOM}};
  bht_120 = _RAND_120[2:0];
  _RAND_121 = {1{`RANDOM}};
  bht_121 = _RAND_121[2:0];
  _RAND_122 = {1{`RANDOM}};
  bht_122 = _RAND_122[2:0];
  _RAND_123 = {1{`RANDOM}};
  bht_123 = _RAND_123[2:0];
  _RAND_124 = {1{`RANDOM}};
  bht_124 = _RAND_124[2:0];
  _RAND_125 = {1{`RANDOM}};
  bht_125 = _RAND_125[2:0];
  _RAND_126 = {1{`RANDOM}};
  bht_126 = _RAND_126[2:0];
  _RAND_127 = {1{`RANDOM}};
  bht_127 = _RAND_127[2:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    bht_0 = 3'h0;
  end
  if (reset) begin
    bht_1 = 3'h0;
  end
  if (reset) begin
    bht_2 = 3'h0;
  end
  if (reset) begin
    bht_3 = 3'h0;
  end
  if (reset) begin
    bht_4 = 3'h0;
  end
  if (reset) begin
    bht_5 = 3'h0;
  end
  if (reset) begin
    bht_6 = 3'h0;
  end
  if (reset) begin
    bht_7 = 3'h0;
  end
  if (reset) begin
    bht_8 = 3'h0;
  end
  if (reset) begin
    bht_9 = 3'h0;
  end
  if (reset) begin
    bht_10 = 3'h0;
  end
  if (reset) begin
    bht_11 = 3'h0;
  end
  if (reset) begin
    bht_12 = 3'h0;
  end
  if (reset) begin
    bht_13 = 3'h0;
  end
  if (reset) begin
    bht_14 = 3'h0;
  end
  if (reset) begin
    bht_15 = 3'h0;
  end
  if (reset) begin
    bht_16 = 3'h0;
  end
  if (reset) begin
    bht_17 = 3'h0;
  end
  if (reset) begin
    bht_18 = 3'h0;
  end
  if (reset) begin
    bht_19 = 3'h0;
  end
  if (reset) begin
    bht_20 = 3'h0;
  end
  if (reset) begin
    bht_21 = 3'h0;
  end
  if (reset) begin
    bht_22 = 3'h0;
  end
  if (reset) begin
    bht_23 = 3'h0;
  end
  if (reset) begin
    bht_24 = 3'h0;
  end
  if (reset) begin
    bht_25 = 3'h0;
  end
  if (reset) begin
    bht_26 = 3'h0;
  end
  if (reset) begin
    bht_27 = 3'h0;
  end
  if (reset) begin
    bht_28 = 3'h0;
  end
  if (reset) begin
    bht_29 = 3'h0;
  end
  if (reset) begin
    bht_30 = 3'h0;
  end
  if (reset) begin
    bht_31 = 3'h0;
  end
  if (reset) begin
    bht_32 = 3'h0;
  end
  if (reset) begin
    bht_33 = 3'h0;
  end
  if (reset) begin
    bht_34 = 3'h0;
  end
  if (reset) begin
    bht_35 = 3'h0;
  end
  if (reset) begin
    bht_36 = 3'h0;
  end
  if (reset) begin
    bht_37 = 3'h0;
  end
  if (reset) begin
    bht_38 = 3'h0;
  end
  if (reset) begin
    bht_39 = 3'h0;
  end
  if (reset) begin
    bht_40 = 3'h0;
  end
  if (reset) begin
    bht_41 = 3'h0;
  end
  if (reset) begin
    bht_42 = 3'h0;
  end
  if (reset) begin
    bht_43 = 3'h0;
  end
  if (reset) begin
    bht_44 = 3'h0;
  end
  if (reset) begin
    bht_45 = 3'h0;
  end
  if (reset) begin
    bht_46 = 3'h0;
  end
  if (reset) begin
    bht_47 = 3'h0;
  end
  if (reset) begin
    bht_48 = 3'h0;
  end
  if (reset) begin
    bht_49 = 3'h0;
  end
  if (reset) begin
    bht_50 = 3'h0;
  end
  if (reset) begin
    bht_51 = 3'h0;
  end
  if (reset) begin
    bht_52 = 3'h0;
  end
  if (reset) begin
    bht_53 = 3'h0;
  end
  if (reset) begin
    bht_54 = 3'h0;
  end
  if (reset) begin
    bht_55 = 3'h0;
  end
  if (reset) begin
    bht_56 = 3'h0;
  end
  if (reset) begin
    bht_57 = 3'h0;
  end
  if (reset) begin
    bht_58 = 3'h0;
  end
  if (reset) begin
    bht_59 = 3'h0;
  end
  if (reset) begin
    bht_60 = 3'h0;
  end
  if (reset) begin
    bht_61 = 3'h0;
  end
  if (reset) begin
    bht_62 = 3'h0;
  end
  if (reset) begin
    bht_63 = 3'h0;
  end
  if (reset) begin
    bht_64 = 3'h0;
  end
  if (reset) begin
    bht_65 = 3'h0;
  end
  if (reset) begin
    bht_66 = 3'h0;
  end
  if (reset) begin
    bht_67 = 3'h0;
  end
  if (reset) begin
    bht_68 = 3'h0;
  end
  if (reset) begin
    bht_69 = 3'h0;
  end
  if (reset) begin
    bht_70 = 3'h0;
  end
  if (reset) begin
    bht_71 = 3'h0;
  end
  if (reset) begin
    bht_72 = 3'h0;
  end
  if (reset) begin
    bht_73 = 3'h0;
  end
  if (reset) begin
    bht_74 = 3'h0;
  end
  if (reset) begin
    bht_75 = 3'h0;
  end
  if (reset) begin
    bht_76 = 3'h0;
  end
  if (reset) begin
    bht_77 = 3'h0;
  end
  if (reset) begin
    bht_78 = 3'h0;
  end
  if (reset) begin
    bht_79 = 3'h0;
  end
  if (reset) begin
    bht_80 = 3'h0;
  end
  if (reset) begin
    bht_81 = 3'h0;
  end
  if (reset) begin
    bht_82 = 3'h0;
  end
  if (reset) begin
    bht_83 = 3'h0;
  end
  if (reset) begin
    bht_84 = 3'h0;
  end
  if (reset) begin
    bht_85 = 3'h0;
  end
  if (reset) begin
    bht_86 = 3'h0;
  end
  if (reset) begin
    bht_87 = 3'h0;
  end
  if (reset) begin
    bht_88 = 3'h0;
  end
  if (reset) begin
    bht_89 = 3'h0;
  end
  if (reset) begin
    bht_90 = 3'h0;
  end
  if (reset) begin
    bht_91 = 3'h0;
  end
  if (reset) begin
    bht_92 = 3'h0;
  end
  if (reset) begin
    bht_93 = 3'h0;
  end
  if (reset) begin
    bht_94 = 3'h0;
  end
  if (reset) begin
    bht_95 = 3'h0;
  end
  if (reset) begin
    bht_96 = 3'h0;
  end
  if (reset) begin
    bht_97 = 3'h0;
  end
  if (reset) begin
    bht_98 = 3'h0;
  end
  if (reset) begin
    bht_99 = 3'h0;
  end
  if (reset) begin
    bht_100 = 3'h0;
  end
  if (reset) begin
    bht_101 = 3'h0;
  end
  if (reset) begin
    bht_102 = 3'h0;
  end
  if (reset) begin
    bht_103 = 3'h0;
  end
  if (reset) begin
    bht_104 = 3'h0;
  end
  if (reset) begin
    bht_105 = 3'h0;
  end
  if (reset) begin
    bht_106 = 3'h0;
  end
  if (reset) begin
    bht_107 = 3'h0;
  end
  if (reset) begin
    bht_108 = 3'h0;
  end
  if (reset) begin
    bht_109 = 3'h0;
  end
  if (reset) begin
    bht_110 = 3'h0;
  end
  if (reset) begin
    bht_111 = 3'h0;
  end
  if (reset) begin
    bht_112 = 3'h0;
  end
  if (reset) begin
    bht_113 = 3'h0;
  end
  if (reset) begin
    bht_114 = 3'h0;
  end
  if (reset) begin
    bht_115 = 3'h0;
  end
  if (reset) begin
    bht_116 = 3'h0;
  end
  if (reset) begin
    bht_117 = 3'h0;
  end
  if (reset) begin
    bht_118 = 3'h0;
  end
  if (reset) begin
    bht_119 = 3'h0;
  end
  if (reset) begin
    bht_120 = 3'h0;
  end
  if (reset) begin
    bht_121 = 3'h0;
  end
  if (reset) begin
    bht_122 = 3'h0;
  end
  if (reset) begin
    bht_123 = 3'h0;
  end
  if (reset) begin
    bht_124 = 3'h0;
  end
  if (reset) begin
    bht_125 = 3'h0;
  end
  if (reset) begin
    bht_126 = 3'h0;
  end
  if (reset) begin
    bht_127 = 3'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BHT_banks_oneissue(
  input        clock,
  input        reset,
  input  [1:0] io_ar_bank_sel,
  input  [6:0] io_ar_addr_L,
  input  [6:0] io_aw_addr,
  input        io_write,
  input  [2:0] io_in,
  output [2:0] io_out_L
);
  wire  BHT_clock; // @[BHT.scala 84:54]
  wire  BHT_reset; // @[BHT.scala 84:54]
  wire [6:0] BHT_io_ar_addr; // @[BHT.scala 84:54]
  wire [6:0] BHT_io_aw_addr; // @[BHT.scala 84:54]
  wire  BHT_io_write; // @[BHT.scala 84:54]
  wire [2:0] BHT_io_in; // @[BHT.scala 84:54]
  wire [2:0] BHT_io_out; // @[BHT.scala 84:54]
  wire  BHT_1_clock; // @[BHT.scala 84:54]
  wire  BHT_1_reset; // @[BHT.scala 84:54]
  wire [6:0] BHT_1_io_ar_addr; // @[BHT.scala 84:54]
  wire [6:0] BHT_1_io_aw_addr; // @[BHT.scala 84:54]
  wire  BHT_1_io_write; // @[BHT.scala 84:54]
  wire [2:0] BHT_1_io_in; // @[BHT.scala 84:54]
  wire [2:0] BHT_1_io_out; // @[BHT.scala 84:54]
  wire  BHT_2_clock; // @[BHT.scala 84:54]
  wire  BHT_2_reset; // @[BHT.scala 84:54]
  wire [6:0] BHT_2_io_ar_addr; // @[BHT.scala 84:54]
  wire [6:0] BHT_2_io_aw_addr; // @[BHT.scala 84:54]
  wire  BHT_2_io_write; // @[BHT.scala 84:54]
  wire [2:0] BHT_2_io_in; // @[BHT.scala 84:54]
  wire [2:0] BHT_2_io_out; // @[BHT.scala 84:54]
  wire  BHT_3_clock; // @[BHT.scala 84:54]
  wire  BHT_3_reset; // @[BHT.scala 84:54]
  wire [6:0] BHT_3_io_ar_addr; // @[BHT.scala 84:54]
  wire [6:0] BHT_3_io_aw_addr; // @[BHT.scala 84:54]
  wire  BHT_3_io_write; // @[BHT.scala 84:54]
  wire [2:0] BHT_3_io_in; // @[BHT.scala 84:54]
  wire [2:0] BHT_3_io_out; // @[BHT.scala 84:54]
  wire [2:0] bht_banks_0_out = BHT_io_out; // @[BHT.scala 84:{28,28}]
  wire [2:0] bht_banks_1_out = BHT_1_io_out; // @[BHT.scala 84:{28,28}]
  wire [2:0] _GEN_1 = 2'h1 == io_ar_bank_sel ? bht_banks_1_out : bht_banks_0_out; // @[BHT.scala 96:{14,14}]
  wire [2:0] bht_banks_2_out = BHT_2_io_out; // @[BHT.scala 84:{28,28}]
  wire [2:0] _GEN_2 = 2'h2 == io_ar_bank_sel ? bht_banks_2_out : _GEN_1; // @[BHT.scala 96:{14,14}]
  wire [2:0] bht_banks_3_out = BHT_3_io_out; // @[BHT.scala 84:{28,28}]
  BHT BHT ( // @[BHT.scala 84:54]
    .clock(BHT_clock),
    .reset(BHT_reset),
    .io_ar_addr(BHT_io_ar_addr),
    .io_aw_addr(BHT_io_aw_addr),
    .io_write(BHT_io_write),
    .io_in(BHT_io_in),
    .io_out(BHT_io_out)
  );
  BHT BHT_1 ( // @[BHT.scala 84:54]
    .clock(BHT_1_clock),
    .reset(BHT_1_reset),
    .io_ar_addr(BHT_1_io_ar_addr),
    .io_aw_addr(BHT_1_io_aw_addr),
    .io_write(BHT_1_io_write),
    .io_in(BHT_1_io_in),
    .io_out(BHT_1_io_out)
  );
  BHT BHT_2 ( // @[BHT.scala 84:54]
    .clock(BHT_2_clock),
    .reset(BHT_2_reset),
    .io_ar_addr(BHT_2_io_ar_addr),
    .io_aw_addr(BHT_2_io_aw_addr),
    .io_write(BHT_2_io_write),
    .io_in(BHT_2_io_in),
    .io_out(BHT_2_io_out)
  );
  BHT BHT_3 ( // @[BHT.scala 84:54]
    .clock(BHT_3_clock),
    .reset(BHT_3_reset),
    .io_ar_addr(BHT_3_io_ar_addr),
    .io_aw_addr(BHT_3_io_aw_addr),
    .io_write(BHT_3_io_write),
    .io_in(BHT_3_io_in),
    .io_out(BHT_3_io_out)
  );
  assign io_out_L = 2'h3 == io_ar_bank_sel ? bht_banks_3_out : _GEN_2; // @[BHT.scala 96:{14,14}]
  assign BHT_clock = clock;
  assign BHT_reset = reset;
  assign BHT_io_ar_addr = io_ar_addr_L; // @[BHT.scala 84:28 88:30]
  assign BHT_io_aw_addr = io_aw_addr; // @[BHT.scala 84:28 94:30]
  assign BHT_io_write = io_ar_bank_sel == 2'h0 & io_write; // @[BHT.scala 86:59]
  assign BHT_io_in = io_in; // @[BHT.scala 84:28 87:25]
  assign BHT_1_clock = clock;
  assign BHT_1_reset = reset;
  assign BHT_1_io_ar_addr = io_ar_addr_L; // @[BHT.scala 84:28 88:30]
  assign BHT_1_io_aw_addr = io_aw_addr; // @[BHT.scala 84:28 94:30]
  assign BHT_1_io_write = io_ar_bank_sel == 2'h1 & io_write; // @[BHT.scala 86:59]
  assign BHT_1_io_in = io_in; // @[BHT.scala 84:28 87:25]
  assign BHT_2_clock = clock;
  assign BHT_2_reset = reset;
  assign BHT_2_io_ar_addr = io_ar_addr_L; // @[BHT.scala 84:28 88:30]
  assign BHT_2_io_aw_addr = io_aw_addr; // @[BHT.scala 84:28 94:30]
  assign BHT_2_io_write = io_ar_bank_sel == 2'h2 & io_write; // @[BHT.scala 86:59]
  assign BHT_2_io_in = io_in; // @[BHT.scala 84:28 87:25]
  assign BHT_3_clock = clock;
  assign BHT_3_reset = reset;
  assign BHT_3_io_ar_addr = io_ar_addr_L; // @[BHT.scala 84:28 88:30]
  assign BHT_3_io_aw_addr = io_aw_addr; // @[BHT.scala 84:28 94:30]
  assign BHT_3_io_write = io_ar_bank_sel == 2'h3 & io_write; // @[BHT.scala 86:59]
  assign BHT_3_io_in = io_in; // @[BHT.scala 84:28 87:25]
endmodule
module Look_up_table_read_first__32(
  input        clock,
  input        reset,
  input  [8:0] io_ar_addr,
  input  [8:0] io_aw_addr,
  input        io_write,
  input  [7:0] io_in,
  output [7:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] btb_0; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_1; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_2; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_3; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_4; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_5; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_6; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_7; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_8; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_9; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_10; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_11; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_12; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_13; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_14; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_15; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_16; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_17; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_18; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_19; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_20; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_21; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_22; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_23; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_24; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_25; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_26; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_27; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_28; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_29; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_30; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_31; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_32; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_33; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_34; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_35; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_36; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_37; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_38; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_39; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_40; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_41; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_42; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_43; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_44; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_45; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_46; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_47; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_48; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_49; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_50; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_51; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_52; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_53; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_54; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_55; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_56; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_57; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_58; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_59; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_60; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_61; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_62; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_63; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_64; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_65; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_66; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_67; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_68; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_69; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_70; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_71; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_72; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_73; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_74; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_75; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_76; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_77; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_78; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_79; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_80; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_81; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_82; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_83; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_84; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_85; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_86; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_87; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_88; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_89; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_90; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_91; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_92; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_93; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_94; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_95; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_96; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_97; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_98; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_99; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_100; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_101; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_102; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_103; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_104; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_105; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_106; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_107; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_108; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_109; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_110; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_111; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_112; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_113; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_114; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_115; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_116; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_117; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_118; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_119; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_120; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_121; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_122; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_123; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_124; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_125; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_126; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_127; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_128; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_129; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_130; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_131; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_132; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_133; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_134; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_135; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_136; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_137; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_138; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_139; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_140; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_141; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_142; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_143; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_144; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_145; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_146; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_147; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_148; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_149; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_150; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_151; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_152; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_153; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_154; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_155; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_156; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_157; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_158; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_159; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_160; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_161; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_162; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_163; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_164; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_165; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_166; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_167; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_168; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_169; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_170; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_171; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_172; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_173; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_174; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_175; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_176; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_177; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_178; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_179; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_180; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_181; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_182; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_183; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_184; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_185; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_186; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_187; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_188; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_189; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_190; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_191; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_192; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_193; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_194; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_195; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_196; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_197; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_198; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_199; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_200; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_201; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_202; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_203; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_204; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_205; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_206; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_207; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_208; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_209; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_210; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_211; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_212; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_213; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_214; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_215; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_216; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_217; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_218; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_219; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_220; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_221; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_222; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_223; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_224; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_225; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_226; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_227; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_228; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_229; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_230; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_231; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_232; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_233; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_234; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_235; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_236; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_237; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_238; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_239; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_240; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_241; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_242; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_243; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_244; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_245; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_246; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_247; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_248; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_249; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_250; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_251; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_252; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_253; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_254; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_255; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_256; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_257; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_258; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_259; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_260; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_261; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_262; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_263; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_264; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_265; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_266; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_267; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_268; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_269; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_270; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_271; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_272; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_273; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_274; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_275; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_276; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_277; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_278; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_279; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_280; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_281; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_282; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_283; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_284; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_285; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_286; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_287; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_288; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_289; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_290; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_291; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_292; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_293; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_294; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_295; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_296; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_297; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_298; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_299; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_300; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_301; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_302; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_303; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_304; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_305; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_306; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_307; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_308; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_309; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_310; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_311; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_312; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_313; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_314; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_315; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_316; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_317; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_318; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_319; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_320; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_321; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_322; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_323; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_324; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_325; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_326; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_327; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_328; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_329; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_330; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_331; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_332; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_333; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_334; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_335; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_336; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_337; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_338; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_339; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_340; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_341; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_342; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_343; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_344; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_345; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_346; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_347; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_348; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_349; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_350; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_351; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_352; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_353; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_354; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_355; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_356; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_357; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_358; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_359; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_360; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_361; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_362; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_363; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_364; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_365; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_366; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_367; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_368; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_369; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_370; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_371; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_372; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_373; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_374; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_375; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_376; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_377; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_378; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_379; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_380; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_381; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_382; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_383; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_384; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_385; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_386; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_387; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_388; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_389; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_390; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_391; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_392; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_393; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_394; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_395; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_396; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_397; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_398; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_399; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_400; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_401; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_402; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_403; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_404; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_405; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_406; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_407; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_408; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_409; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_410; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_411; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_412; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_413; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_414; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_415; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_416; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_417; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_418; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_419; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_420; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_421; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_422; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_423; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_424; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_425; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_426; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_427; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_428; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_429; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_430; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_431; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_432; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_433; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_434; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_435; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_436; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_437; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_438; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_439; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_440; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_441; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_442; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_443; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_444; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_445; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_446; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_447; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_448; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_449; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_450; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_451; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_452; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_453; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_454; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_455; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_456; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_457; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_458; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_459; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_460; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_461; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_462; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_463; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_464; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_465; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_466; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_467; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_468; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_469; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_470; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_471; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_472; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_473; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_474; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_475; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_476; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_477; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_478; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_479; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_480; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_481; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_482; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_483; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_484; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_485; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_486; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_487; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_488; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_489; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_490; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_491; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_492; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_493; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_494; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_495; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_496; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_497; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_498; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_499; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_500; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_501; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_502; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_503; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_504; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_505; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_506; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_507; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_508; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_509; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_510; // @[ports_lookup_table.scala 81:22]
  reg [7:0] btb_511; // @[ports_lookup_table.scala 81:22]
  wire [7:0] _GEN_1 = 9'h1 == io_ar_addr ? btb_1 : btb_0; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_2 = 9'h2 == io_ar_addr ? btb_2 : _GEN_1; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_3 = 9'h3 == io_ar_addr ? btb_3 : _GEN_2; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_4 = 9'h4 == io_ar_addr ? btb_4 : _GEN_3; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_5 = 9'h5 == io_ar_addr ? btb_5 : _GEN_4; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_6 = 9'h6 == io_ar_addr ? btb_6 : _GEN_5; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_7 = 9'h7 == io_ar_addr ? btb_7 : _GEN_6; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_8 = 9'h8 == io_ar_addr ? btb_8 : _GEN_7; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_9 = 9'h9 == io_ar_addr ? btb_9 : _GEN_8; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_10 = 9'ha == io_ar_addr ? btb_10 : _GEN_9; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_11 = 9'hb == io_ar_addr ? btb_11 : _GEN_10; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_12 = 9'hc == io_ar_addr ? btb_12 : _GEN_11; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_13 = 9'hd == io_ar_addr ? btb_13 : _GEN_12; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_14 = 9'he == io_ar_addr ? btb_14 : _GEN_13; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_15 = 9'hf == io_ar_addr ? btb_15 : _GEN_14; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_16 = 9'h10 == io_ar_addr ? btb_16 : _GEN_15; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_17 = 9'h11 == io_ar_addr ? btb_17 : _GEN_16; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_18 = 9'h12 == io_ar_addr ? btb_18 : _GEN_17; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_19 = 9'h13 == io_ar_addr ? btb_19 : _GEN_18; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_20 = 9'h14 == io_ar_addr ? btb_20 : _GEN_19; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_21 = 9'h15 == io_ar_addr ? btb_21 : _GEN_20; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_22 = 9'h16 == io_ar_addr ? btb_22 : _GEN_21; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_23 = 9'h17 == io_ar_addr ? btb_23 : _GEN_22; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_24 = 9'h18 == io_ar_addr ? btb_24 : _GEN_23; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_25 = 9'h19 == io_ar_addr ? btb_25 : _GEN_24; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_26 = 9'h1a == io_ar_addr ? btb_26 : _GEN_25; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_27 = 9'h1b == io_ar_addr ? btb_27 : _GEN_26; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_28 = 9'h1c == io_ar_addr ? btb_28 : _GEN_27; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_29 = 9'h1d == io_ar_addr ? btb_29 : _GEN_28; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_30 = 9'h1e == io_ar_addr ? btb_30 : _GEN_29; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_31 = 9'h1f == io_ar_addr ? btb_31 : _GEN_30; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_32 = 9'h20 == io_ar_addr ? btb_32 : _GEN_31; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_33 = 9'h21 == io_ar_addr ? btb_33 : _GEN_32; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_34 = 9'h22 == io_ar_addr ? btb_34 : _GEN_33; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_35 = 9'h23 == io_ar_addr ? btb_35 : _GEN_34; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_36 = 9'h24 == io_ar_addr ? btb_36 : _GEN_35; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_37 = 9'h25 == io_ar_addr ? btb_37 : _GEN_36; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_38 = 9'h26 == io_ar_addr ? btb_38 : _GEN_37; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_39 = 9'h27 == io_ar_addr ? btb_39 : _GEN_38; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_40 = 9'h28 == io_ar_addr ? btb_40 : _GEN_39; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_41 = 9'h29 == io_ar_addr ? btb_41 : _GEN_40; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_42 = 9'h2a == io_ar_addr ? btb_42 : _GEN_41; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_43 = 9'h2b == io_ar_addr ? btb_43 : _GEN_42; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_44 = 9'h2c == io_ar_addr ? btb_44 : _GEN_43; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_45 = 9'h2d == io_ar_addr ? btb_45 : _GEN_44; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_46 = 9'h2e == io_ar_addr ? btb_46 : _GEN_45; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_47 = 9'h2f == io_ar_addr ? btb_47 : _GEN_46; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_48 = 9'h30 == io_ar_addr ? btb_48 : _GEN_47; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_49 = 9'h31 == io_ar_addr ? btb_49 : _GEN_48; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_50 = 9'h32 == io_ar_addr ? btb_50 : _GEN_49; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_51 = 9'h33 == io_ar_addr ? btb_51 : _GEN_50; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_52 = 9'h34 == io_ar_addr ? btb_52 : _GEN_51; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_53 = 9'h35 == io_ar_addr ? btb_53 : _GEN_52; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_54 = 9'h36 == io_ar_addr ? btb_54 : _GEN_53; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_55 = 9'h37 == io_ar_addr ? btb_55 : _GEN_54; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_56 = 9'h38 == io_ar_addr ? btb_56 : _GEN_55; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_57 = 9'h39 == io_ar_addr ? btb_57 : _GEN_56; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_58 = 9'h3a == io_ar_addr ? btb_58 : _GEN_57; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_59 = 9'h3b == io_ar_addr ? btb_59 : _GEN_58; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_60 = 9'h3c == io_ar_addr ? btb_60 : _GEN_59; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_61 = 9'h3d == io_ar_addr ? btb_61 : _GEN_60; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_62 = 9'h3e == io_ar_addr ? btb_62 : _GEN_61; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_63 = 9'h3f == io_ar_addr ? btb_63 : _GEN_62; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_64 = 9'h40 == io_ar_addr ? btb_64 : _GEN_63; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_65 = 9'h41 == io_ar_addr ? btb_65 : _GEN_64; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_66 = 9'h42 == io_ar_addr ? btb_66 : _GEN_65; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_67 = 9'h43 == io_ar_addr ? btb_67 : _GEN_66; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_68 = 9'h44 == io_ar_addr ? btb_68 : _GEN_67; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_69 = 9'h45 == io_ar_addr ? btb_69 : _GEN_68; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_70 = 9'h46 == io_ar_addr ? btb_70 : _GEN_69; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_71 = 9'h47 == io_ar_addr ? btb_71 : _GEN_70; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_72 = 9'h48 == io_ar_addr ? btb_72 : _GEN_71; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_73 = 9'h49 == io_ar_addr ? btb_73 : _GEN_72; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_74 = 9'h4a == io_ar_addr ? btb_74 : _GEN_73; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_75 = 9'h4b == io_ar_addr ? btb_75 : _GEN_74; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_76 = 9'h4c == io_ar_addr ? btb_76 : _GEN_75; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_77 = 9'h4d == io_ar_addr ? btb_77 : _GEN_76; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_78 = 9'h4e == io_ar_addr ? btb_78 : _GEN_77; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_79 = 9'h4f == io_ar_addr ? btb_79 : _GEN_78; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_80 = 9'h50 == io_ar_addr ? btb_80 : _GEN_79; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_81 = 9'h51 == io_ar_addr ? btb_81 : _GEN_80; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_82 = 9'h52 == io_ar_addr ? btb_82 : _GEN_81; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_83 = 9'h53 == io_ar_addr ? btb_83 : _GEN_82; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_84 = 9'h54 == io_ar_addr ? btb_84 : _GEN_83; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_85 = 9'h55 == io_ar_addr ? btb_85 : _GEN_84; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_86 = 9'h56 == io_ar_addr ? btb_86 : _GEN_85; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_87 = 9'h57 == io_ar_addr ? btb_87 : _GEN_86; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_88 = 9'h58 == io_ar_addr ? btb_88 : _GEN_87; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_89 = 9'h59 == io_ar_addr ? btb_89 : _GEN_88; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_90 = 9'h5a == io_ar_addr ? btb_90 : _GEN_89; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_91 = 9'h5b == io_ar_addr ? btb_91 : _GEN_90; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_92 = 9'h5c == io_ar_addr ? btb_92 : _GEN_91; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_93 = 9'h5d == io_ar_addr ? btb_93 : _GEN_92; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_94 = 9'h5e == io_ar_addr ? btb_94 : _GEN_93; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_95 = 9'h5f == io_ar_addr ? btb_95 : _GEN_94; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_96 = 9'h60 == io_ar_addr ? btb_96 : _GEN_95; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_97 = 9'h61 == io_ar_addr ? btb_97 : _GEN_96; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_98 = 9'h62 == io_ar_addr ? btb_98 : _GEN_97; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_99 = 9'h63 == io_ar_addr ? btb_99 : _GEN_98; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_100 = 9'h64 == io_ar_addr ? btb_100 : _GEN_99; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_101 = 9'h65 == io_ar_addr ? btb_101 : _GEN_100; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_102 = 9'h66 == io_ar_addr ? btb_102 : _GEN_101; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_103 = 9'h67 == io_ar_addr ? btb_103 : _GEN_102; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_104 = 9'h68 == io_ar_addr ? btb_104 : _GEN_103; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_105 = 9'h69 == io_ar_addr ? btb_105 : _GEN_104; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_106 = 9'h6a == io_ar_addr ? btb_106 : _GEN_105; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_107 = 9'h6b == io_ar_addr ? btb_107 : _GEN_106; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_108 = 9'h6c == io_ar_addr ? btb_108 : _GEN_107; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_109 = 9'h6d == io_ar_addr ? btb_109 : _GEN_108; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_110 = 9'h6e == io_ar_addr ? btb_110 : _GEN_109; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_111 = 9'h6f == io_ar_addr ? btb_111 : _GEN_110; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_112 = 9'h70 == io_ar_addr ? btb_112 : _GEN_111; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_113 = 9'h71 == io_ar_addr ? btb_113 : _GEN_112; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_114 = 9'h72 == io_ar_addr ? btb_114 : _GEN_113; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_115 = 9'h73 == io_ar_addr ? btb_115 : _GEN_114; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_116 = 9'h74 == io_ar_addr ? btb_116 : _GEN_115; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_117 = 9'h75 == io_ar_addr ? btb_117 : _GEN_116; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_118 = 9'h76 == io_ar_addr ? btb_118 : _GEN_117; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_119 = 9'h77 == io_ar_addr ? btb_119 : _GEN_118; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_120 = 9'h78 == io_ar_addr ? btb_120 : _GEN_119; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_121 = 9'h79 == io_ar_addr ? btb_121 : _GEN_120; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_122 = 9'h7a == io_ar_addr ? btb_122 : _GEN_121; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_123 = 9'h7b == io_ar_addr ? btb_123 : _GEN_122; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_124 = 9'h7c == io_ar_addr ? btb_124 : _GEN_123; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_125 = 9'h7d == io_ar_addr ? btb_125 : _GEN_124; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_126 = 9'h7e == io_ar_addr ? btb_126 : _GEN_125; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_127 = 9'h7f == io_ar_addr ? btb_127 : _GEN_126; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_128 = 9'h80 == io_ar_addr ? btb_128 : _GEN_127; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_129 = 9'h81 == io_ar_addr ? btb_129 : _GEN_128; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_130 = 9'h82 == io_ar_addr ? btb_130 : _GEN_129; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_131 = 9'h83 == io_ar_addr ? btb_131 : _GEN_130; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_132 = 9'h84 == io_ar_addr ? btb_132 : _GEN_131; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_133 = 9'h85 == io_ar_addr ? btb_133 : _GEN_132; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_134 = 9'h86 == io_ar_addr ? btb_134 : _GEN_133; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_135 = 9'h87 == io_ar_addr ? btb_135 : _GEN_134; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_136 = 9'h88 == io_ar_addr ? btb_136 : _GEN_135; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_137 = 9'h89 == io_ar_addr ? btb_137 : _GEN_136; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_138 = 9'h8a == io_ar_addr ? btb_138 : _GEN_137; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_139 = 9'h8b == io_ar_addr ? btb_139 : _GEN_138; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_140 = 9'h8c == io_ar_addr ? btb_140 : _GEN_139; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_141 = 9'h8d == io_ar_addr ? btb_141 : _GEN_140; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_142 = 9'h8e == io_ar_addr ? btb_142 : _GEN_141; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_143 = 9'h8f == io_ar_addr ? btb_143 : _GEN_142; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_144 = 9'h90 == io_ar_addr ? btb_144 : _GEN_143; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_145 = 9'h91 == io_ar_addr ? btb_145 : _GEN_144; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_146 = 9'h92 == io_ar_addr ? btb_146 : _GEN_145; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_147 = 9'h93 == io_ar_addr ? btb_147 : _GEN_146; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_148 = 9'h94 == io_ar_addr ? btb_148 : _GEN_147; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_149 = 9'h95 == io_ar_addr ? btb_149 : _GEN_148; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_150 = 9'h96 == io_ar_addr ? btb_150 : _GEN_149; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_151 = 9'h97 == io_ar_addr ? btb_151 : _GEN_150; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_152 = 9'h98 == io_ar_addr ? btb_152 : _GEN_151; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_153 = 9'h99 == io_ar_addr ? btb_153 : _GEN_152; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_154 = 9'h9a == io_ar_addr ? btb_154 : _GEN_153; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_155 = 9'h9b == io_ar_addr ? btb_155 : _GEN_154; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_156 = 9'h9c == io_ar_addr ? btb_156 : _GEN_155; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_157 = 9'h9d == io_ar_addr ? btb_157 : _GEN_156; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_158 = 9'h9e == io_ar_addr ? btb_158 : _GEN_157; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_159 = 9'h9f == io_ar_addr ? btb_159 : _GEN_158; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_160 = 9'ha0 == io_ar_addr ? btb_160 : _GEN_159; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_161 = 9'ha1 == io_ar_addr ? btb_161 : _GEN_160; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_162 = 9'ha2 == io_ar_addr ? btb_162 : _GEN_161; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_163 = 9'ha3 == io_ar_addr ? btb_163 : _GEN_162; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_164 = 9'ha4 == io_ar_addr ? btb_164 : _GEN_163; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_165 = 9'ha5 == io_ar_addr ? btb_165 : _GEN_164; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_166 = 9'ha6 == io_ar_addr ? btb_166 : _GEN_165; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_167 = 9'ha7 == io_ar_addr ? btb_167 : _GEN_166; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_168 = 9'ha8 == io_ar_addr ? btb_168 : _GEN_167; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_169 = 9'ha9 == io_ar_addr ? btb_169 : _GEN_168; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_170 = 9'haa == io_ar_addr ? btb_170 : _GEN_169; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_171 = 9'hab == io_ar_addr ? btb_171 : _GEN_170; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_172 = 9'hac == io_ar_addr ? btb_172 : _GEN_171; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_173 = 9'had == io_ar_addr ? btb_173 : _GEN_172; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_174 = 9'hae == io_ar_addr ? btb_174 : _GEN_173; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_175 = 9'haf == io_ar_addr ? btb_175 : _GEN_174; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_176 = 9'hb0 == io_ar_addr ? btb_176 : _GEN_175; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_177 = 9'hb1 == io_ar_addr ? btb_177 : _GEN_176; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_178 = 9'hb2 == io_ar_addr ? btb_178 : _GEN_177; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_179 = 9'hb3 == io_ar_addr ? btb_179 : _GEN_178; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_180 = 9'hb4 == io_ar_addr ? btb_180 : _GEN_179; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_181 = 9'hb5 == io_ar_addr ? btb_181 : _GEN_180; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_182 = 9'hb6 == io_ar_addr ? btb_182 : _GEN_181; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_183 = 9'hb7 == io_ar_addr ? btb_183 : _GEN_182; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_184 = 9'hb8 == io_ar_addr ? btb_184 : _GEN_183; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_185 = 9'hb9 == io_ar_addr ? btb_185 : _GEN_184; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_186 = 9'hba == io_ar_addr ? btb_186 : _GEN_185; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_187 = 9'hbb == io_ar_addr ? btb_187 : _GEN_186; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_188 = 9'hbc == io_ar_addr ? btb_188 : _GEN_187; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_189 = 9'hbd == io_ar_addr ? btb_189 : _GEN_188; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_190 = 9'hbe == io_ar_addr ? btb_190 : _GEN_189; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_191 = 9'hbf == io_ar_addr ? btb_191 : _GEN_190; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_192 = 9'hc0 == io_ar_addr ? btb_192 : _GEN_191; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_193 = 9'hc1 == io_ar_addr ? btb_193 : _GEN_192; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_194 = 9'hc2 == io_ar_addr ? btb_194 : _GEN_193; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_195 = 9'hc3 == io_ar_addr ? btb_195 : _GEN_194; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_196 = 9'hc4 == io_ar_addr ? btb_196 : _GEN_195; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_197 = 9'hc5 == io_ar_addr ? btb_197 : _GEN_196; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_198 = 9'hc6 == io_ar_addr ? btb_198 : _GEN_197; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_199 = 9'hc7 == io_ar_addr ? btb_199 : _GEN_198; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_200 = 9'hc8 == io_ar_addr ? btb_200 : _GEN_199; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_201 = 9'hc9 == io_ar_addr ? btb_201 : _GEN_200; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_202 = 9'hca == io_ar_addr ? btb_202 : _GEN_201; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_203 = 9'hcb == io_ar_addr ? btb_203 : _GEN_202; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_204 = 9'hcc == io_ar_addr ? btb_204 : _GEN_203; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_205 = 9'hcd == io_ar_addr ? btb_205 : _GEN_204; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_206 = 9'hce == io_ar_addr ? btb_206 : _GEN_205; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_207 = 9'hcf == io_ar_addr ? btb_207 : _GEN_206; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_208 = 9'hd0 == io_ar_addr ? btb_208 : _GEN_207; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_209 = 9'hd1 == io_ar_addr ? btb_209 : _GEN_208; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_210 = 9'hd2 == io_ar_addr ? btb_210 : _GEN_209; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_211 = 9'hd3 == io_ar_addr ? btb_211 : _GEN_210; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_212 = 9'hd4 == io_ar_addr ? btb_212 : _GEN_211; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_213 = 9'hd5 == io_ar_addr ? btb_213 : _GEN_212; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_214 = 9'hd6 == io_ar_addr ? btb_214 : _GEN_213; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_215 = 9'hd7 == io_ar_addr ? btb_215 : _GEN_214; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_216 = 9'hd8 == io_ar_addr ? btb_216 : _GEN_215; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_217 = 9'hd9 == io_ar_addr ? btb_217 : _GEN_216; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_218 = 9'hda == io_ar_addr ? btb_218 : _GEN_217; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_219 = 9'hdb == io_ar_addr ? btb_219 : _GEN_218; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_220 = 9'hdc == io_ar_addr ? btb_220 : _GEN_219; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_221 = 9'hdd == io_ar_addr ? btb_221 : _GEN_220; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_222 = 9'hde == io_ar_addr ? btb_222 : _GEN_221; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_223 = 9'hdf == io_ar_addr ? btb_223 : _GEN_222; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_224 = 9'he0 == io_ar_addr ? btb_224 : _GEN_223; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_225 = 9'he1 == io_ar_addr ? btb_225 : _GEN_224; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_226 = 9'he2 == io_ar_addr ? btb_226 : _GEN_225; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_227 = 9'he3 == io_ar_addr ? btb_227 : _GEN_226; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_228 = 9'he4 == io_ar_addr ? btb_228 : _GEN_227; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_229 = 9'he5 == io_ar_addr ? btb_229 : _GEN_228; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_230 = 9'he6 == io_ar_addr ? btb_230 : _GEN_229; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_231 = 9'he7 == io_ar_addr ? btb_231 : _GEN_230; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_232 = 9'he8 == io_ar_addr ? btb_232 : _GEN_231; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_233 = 9'he9 == io_ar_addr ? btb_233 : _GEN_232; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_234 = 9'hea == io_ar_addr ? btb_234 : _GEN_233; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_235 = 9'heb == io_ar_addr ? btb_235 : _GEN_234; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_236 = 9'hec == io_ar_addr ? btb_236 : _GEN_235; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_237 = 9'hed == io_ar_addr ? btb_237 : _GEN_236; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_238 = 9'hee == io_ar_addr ? btb_238 : _GEN_237; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_239 = 9'hef == io_ar_addr ? btb_239 : _GEN_238; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_240 = 9'hf0 == io_ar_addr ? btb_240 : _GEN_239; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_241 = 9'hf1 == io_ar_addr ? btb_241 : _GEN_240; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_242 = 9'hf2 == io_ar_addr ? btb_242 : _GEN_241; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_243 = 9'hf3 == io_ar_addr ? btb_243 : _GEN_242; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_244 = 9'hf4 == io_ar_addr ? btb_244 : _GEN_243; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_245 = 9'hf5 == io_ar_addr ? btb_245 : _GEN_244; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_246 = 9'hf6 == io_ar_addr ? btb_246 : _GEN_245; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_247 = 9'hf7 == io_ar_addr ? btb_247 : _GEN_246; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_248 = 9'hf8 == io_ar_addr ? btb_248 : _GEN_247; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_249 = 9'hf9 == io_ar_addr ? btb_249 : _GEN_248; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_250 = 9'hfa == io_ar_addr ? btb_250 : _GEN_249; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_251 = 9'hfb == io_ar_addr ? btb_251 : _GEN_250; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_252 = 9'hfc == io_ar_addr ? btb_252 : _GEN_251; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_253 = 9'hfd == io_ar_addr ? btb_253 : _GEN_252; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_254 = 9'hfe == io_ar_addr ? btb_254 : _GEN_253; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_255 = 9'hff == io_ar_addr ? btb_255 : _GEN_254; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_256 = 9'h100 == io_ar_addr ? btb_256 : _GEN_255; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_257 = 9'h101 == io_ar_addr ? btb_257 : _GEN_256; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_258 = 9'h102 == io_ar_addr ? btb_258 : _GEN_257; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_259 = 9'h103 == io_ar_addr ? btb_259 : _GEN_258; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_260 = 9'h104 == io_ar_addr ? btb_260 : _GEN_259; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_261 = 9'h105 == io_ar_addr ? btb_261 : _GEN_260; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_262 = 9'h106 == io_ar_addr ? btb_262 : _GEN_261; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_263 = 9'h107 == io_ar_addr ? btb_263 : _GEN_262; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_264 = 9'h108 == io_ar_addr ? btb_264 : _GEN_263; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_265 = 9'h109 == io_ar_addr ? btb_265 : _GEN_264; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_266 = 9'h10a == io_ar_addr ? btb_266 : _GEN_265; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_267 = 9'h10b == io_ar_addr ? btb_267 : _GEN_266; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_268 = 9'h10c == io_ar_addr ? btb_268 : _GEN_267; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_269 = 9'h10d == io_ar_addr ? btb_269 : _GEN_268; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_270 = 9'h10e == io_ar_addr ? btb_270 : _GEN_269; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_271 = 9'h10f == io_ar_addr ? btb_271 : _GEN_270; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_272 = 9'h110 == io_ar_addr ? btb_272 : _GEN_271; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_273 = 9'h111 == io_ar_addr ? btb_273 : _GEN_272; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_274 = 9'h112 == io_ar_addr ? btb_274 : _GEN_273; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_275 = 9'h113 == io_ar_addr ? btb_275 : _GEN_274; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_276 = 9'h114 == io_ar_addr ? btb_276 : _GEN_275; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_277 = 9'h115 == io_ar_addr ? btb_277 : _GEN_276; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_278 = 9'h116 == io_ar_addr ? btb_278 : _GEN_277; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_279 = 9'h117 == io_ar_addr ? btb_279 : _GEN_278; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_280 = 9'h118 == io_ar_addr ? btb_280 : _GEN_279; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_281 = 9'h119 == io_ar_addr ? btb_281 : _GEN_280; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_282 = 9'h11a == io_ar_addr ? btb_282 : _GEN_281; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_283 = 9'h11b == io_ar_addr ? btb_283 : _GEN_282; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_284 = 9'h11c == io_ar_addr ? btb_284 : _GEN_283; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_285 = 9'h11d == io_ar_addr ? btb_285 : _GEN_284; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_286 = 9'h11e == io_ar_addr ? btb_286 : _GEN_285; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_287 = 9'h11f == io_ar_addr ? btb_287 : _GEN_286; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_288 = 9'h120 == io_ar_addr ? btb_288 : _GEN_287; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_289 = 9'h121 == io_ar_addr ? btb_289 : _GEN_288; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_290 = 9'h122 == io_ar_addr ? btb_290 : _GEN_289; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_291 = 9'h123 == io_ar_addr ? btb_291 : _GEN_290; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_292 = 9'h124 == io_ar_addr ? btb_292 : _GEN_291; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_293 = 9'h125 == io_ar_addr ? btb_293 : _GEN_292; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_294 = 9'h126 == io_ar_addr ? btb_294 : _GEN_293; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_295 = 9'h127 == io_ar_addr ? btb_295 : _GEN_294; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_296 = 9'h128 == io_ar_addr ? btb_296 : _GEN_295; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_297 = 9'h129 == io_ar_addr ? btb_297 : _GEN_296; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_298 = 9'h12a == io_ar_addr ? btb_298 : _GEN_297; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_299 = 9'h12b == io_ar_addr ? btb_299 : _GEN_298; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_300 = 9'h12c == io_ar_addr ? btb_300 : _GEN_299; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_301 = 9'h12d == io_ar_addr ? btb_301 : _GEN_300; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_302 = 9'h12e == io_ar_addr ? btb_302 : _GEN_301; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_303 = 9'h12f == io_ar_addr ? btb_303 : _GEN_302; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_304 = 9'h130 == io_ar_addr ? btb_304 : _GEN_303; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_305 = 9'h131 == io_ar_addr ? btb_305 : _GEN_304; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_306 = 9'h132 == io_ar_addr ? btb_306 : _GEN_305; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_307 = 9'h133 == io_ar_addr ? btb_307 : _GEN_306; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_308 = 9'h134 == io_ar_addr ? btb_308 : _GEN_307; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_309 = 9'h135 == io_ar_addr ? btb_309 : _GEN_308; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_310 = 9'h136 == io_ar_addr ? btb_310 : _GEN_309; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_311 = 9'h137 == io_ar_addr ? btb_311 : _GEN_310; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_312 = 9'h138 == io_ar_addr ? btb_312 : _GEN_311; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_313 = 9'h139 == io_ar_addr ? btb_313 : _GEN_312; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_314 = 9'h13a == io_ar_addr ? btb_314 : _GEN_313; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_315 = 9'h13b == io_ar_addr ? btb_315 : _GEN_314; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_316 = 9'h13c == io_ar_addr ? btb_316 : _GEN_315; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_317 = 9'h13d == io_ar_addr ? btb_317 : _GEN_316; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_318 = 9'h13e == io_ar_addr ? btb_318 : _GEN_317; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_319 = 9'h13f == io_ar_addr ? btb_319 : _GEN_318; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_320 = 9'h140 == io_ar_addr ? btb_320 : _GEN_319; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_321 = 9'h141 == io_ar_addr ? btb_321 : _GEN_320; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_322 = 9'h142 == io_ar_addr ? btb_322 : _GEN_321; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_323 = 9'h143 == io_ar_addr ? btb_323 : _GEN_322; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_324 = 9'h144 == io_ar_addr ? btb_324 : _GEN_323; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_325 = 9'h145 == io_ar_addr ? btb_325 : _GEN_324; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_326 = 9'h146 == io_ar_addr ? btb_326 : _GEN_325; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_327 = 9'h147 == io_ar_addr ? btb_327 : _GEN_326; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_328 = 9'h148 == io_ar_addr ? btb_328 : _GEN_327; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_329 = 9'h149 == io_ar_addr ? btb_329 : _GEN_328; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_330 = 9'h14a == io_ar_addr ? btb_330 : _GEN_329; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_331 = 9'h14b == io_ar_addr ? btb_331 : _GEN_330; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_332 = 9'h14c == io_ar_addr ? btb_332 : _GEN_331; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_333 = 9'h14d == io_ar_addr ? btb_333 : _GEN_332; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_334 = 9'h14e == io_ar_addr ? btb_334 : _GEN_333; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_335 = 9'h14f == io_ar_addr ? btb_335 : _GEN_334; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_336 = 9'h150 == io_ar_addr ? btb_336 : _GEN_335; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_337 = 9'h151 == io_ar_addr ? btb_337 : _GEN_336; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_338 = 9'h152 == io_ar_addr ? btb_338 : _GEN_337; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_339 = 9'h153 == io_ar_addr ? btb_339 : _GEN_338; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_340 = 9'h154 == io_ar_addr ? btb_340 : _GEN_339; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_341 = 9'h155 == io_ar_addr ? btb_341 : _GEN_340; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_342 = 9'h156 == io_ar_addr ? btb_342 : _GEN_341; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_343 = 9'h157 == io_ar_addr ? btb_343 : _GEN_342; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_344 = 9'h158 == io_ar_addr ? btb_344 : _GEN_343; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_345 = 9'h159 == io_ar_addr ? btb_345 : _GEN_344; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_346 = 9'h15a == io_ar_addr ? btb_346 : _GEN_345; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_347 = 9'h15b == io_ar_addr ? btb_347 : _GEN_346; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_348 = 9'h15c == io_ar_addr ? btb_348 : _GEN_347; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_349 = 9'h15d == io_ar_addr ? btb_349 : _GEN_348; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_350 = 9'h15e == io_ar_addr ? btb_350 : _GEN_349; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_351 = 9'h15f == io_ar_addr ? btb_351 : _GEN_350; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_352 = 9'h160 == io_ar_addr ? btb_352 : _GEN_351; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_353 = 9'h161 == io_ar_addr ? btb_353 : _GEN_352; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_354 = 9'h162 == io_ar_addr ? btb_354 : _GEN_353; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_355 = 9'h163 == io_ar_addr ? btb_355 : _GEN_354; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_356 = 9'h164 == io_ar_addr ? btb_356 : _GEN_355; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_357 = 9'h165 == io_ar_addr ? btb_357 : _GEN_356; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_358 = 9'h166 == io_ar_addr ? btb_358 : _GEN_357; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_359 = 9'h167 == io_ar_addr ? btb_359 : _GEN_358; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_360 = 9'h168 == io_ar_addr ? btb_360 : _GEN_359; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_361 = 9'h169 == io_ar_addr ? btb_361 : _GEN_360; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_362 = 9'h16a == io_ar_addr ? btb_362 : _GEN_361; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_363 = 9'h16b == io_ar_addr ? btb_363 : _GEN_362; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_364 = 9'h16c == io_ar_addr ? btb_364 : _GEN_363; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_365 = 9'h16d == io_ar_addr ? btb_365 : _GEN_364; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_366 = 9'h16e == io_ar_addr ? btb_366 : _GEN_365; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_367 = 9'h16f == io_ar_addr ? btb_367 : _GEN_366; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_368 = 9'h170 == io_ar_addr ? btb_368 : _GEN_367; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_369 = 9'h171 == io_ar_addr ? btb_369 : _GEN_368; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_370 = 9'h172 == io_ar_addr ? btb_370 : _GEN_369; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_371 = 9'h173 == io_ar_addr ? btb_371 : _GEN_370; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_372 = 9'h174 == io_ar_addr ? btb_372 : _GEN_371; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_373 = 9'h175 == io_ar_addr ? btb_373 : _GEN_372; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_374 = 9'h176 == io_ar_addr ? btb_374 : _GEN_373; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_375 = 9'h177 == io_ar_addr ? btb_375 : _GEN_374; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_376 = 9'h178 == io_ar_addr ? btb_376 : _GEN_375; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_377 = 9'h179 == io_ar_addr ? btb_377 : _GEN_376; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_378 = 9'h17a == io_ar_addr ? btb_378 : _GEN_377; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_379 = 9'h17b == io_ar_addr ? btb_379 : _GEN_378; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_380 = 9'h17c == io_ar_addr ? btb_380 : _GEN_379; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_381 = 9'h17d == io_ar_addr ? btb_381 : _GEN_380; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_382 = 9'h17e == io_ar_addr ? btb_382 : _GEN_381; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_383 = 9'h17f == io_ar_addr ? btb_383 : _GEN_382; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_384 = 9'h180 == io_ar_addr ? btb_384 : _GEN_383; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_385 = 9'h181 == io_ar_addr ? btb_385 : _GEN_384; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_386 = 9'h182 == io_ar_addr ? btb_386 : _GEN_385; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_387 = 9'h183 == io_ar_addr ? btb_387 : _GEN_386; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_388 = 9'h184 == io_ar_addr ? btb_388 : _GEN_387; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_389 = 9'h185 == io_ar_addr ? btb_389 : _GEN_388; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_390 = 9'h186 == io_ar_addr ? btb_390 : _GEN_389; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_391 = 9'h187 == io_ar_addr ? btb_391 : _GEN_390; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_392 = 9'h188 == io_ar_addr ? btb_392 : _GEN_391; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_393 = 9'h189 == io_ar_addr ? btb_393 : _GEN_392; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_394 = 9'h18a == io_ar_addr ? btb_394 : _GEN_393; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_395 = 9'h18b == io_ar_addr ? btb_395 : _GEN_394; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_396 = 9'h18c == io_ar_addr ? btb_396 : _GEN_395; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_397 = 9'h18d == io_ar_addr ? btb_397 : _GEN_396; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_398 = 9'h18e == io_ar_addr ? btb_398 : _GEN_397; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_399 = 9'h18f == io_ar_addr ? btb_399 : _GEN_398; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_400 = 9'h190 == io_ar_addr ? btb_400 : _GEN_399; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_401 = 9'h191 == io_ar_addr ? btb_401 : _GEN_400; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_402 = 9'h192 == io_ar_addr ? btb_402 : _GEN_401; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_403 = 9'h193 == io_ar_addr ? btb_403 : _GEN_402; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_404 = 9'h194 == io_ar_addr ? btb_404 : _GEN_403; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_405 = 9'h195 == io_ar_addr ? btb_405 : _GEN_404; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_406 = 9'h196 == io_ar_addr ? btb_406 : _GEN_405; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_407 = 9'h197 == io_ar_addr ? btb_407 : _GEN_406; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_408 = 9'h198 == io_ar_addr ? btb_408 : _GEN_407; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_409 = 9'h199 == io_ar_addr ? btb_409 : _GEN_408; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_410 = 9'h19a == io_ar_addr ? btb_410 : _GEN_409; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_411 = 9'h19b == io_ar_addr ? btb_411 : _GEN_410; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_412 = 9'h19c == io_ar_addr ? btb_412 : _GEN_411; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_413 = 9'h19d == io_ar_addr ? btb_413 : _GEN_412; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_414 = 9'h19e == io_ar_addr ? btb_414 : _GEN_413; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_415 = 9'h19f == io_ar_addr ? btb_415 : _GEN_414; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_416 = 9'h1a0 == io_ar_addr ? btb_416 : _GEN_415; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_417 = 9'h1a1 == io_ar_addr ? btb_417 : _GEN_416; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_418 = 9'h1a2 == io_ar_addr ? btb_418 : _GEN_417; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_419 = 9'h1a3 == io_ar_addr ? btb_419 : _GEN_418; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_420 = 9'h1a4 == io_ar_addr ? btb_420 : _GEN_419; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_421 = 9'h1a5 == io_ar_addr ? btb_421 : _GEN_420; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_422 = 9'h1a6 == io_ar_addr ? btb_422 : _GEN_421; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_423 = 9'h1a7 == io_ar_addr ? btb_423 : _GEN_422; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_424 = 9'h1a8 == io_ar_addr ? btb_424 : _GEN_423; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_425 = 9'h1a9 == io_ar_addr ? btb_425 : _GEN_424; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_426 = 9'h1aa == io_ar_addr ? btb_426 : _GEN_425; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_427 = 9'h1ab == io_ar_addr ? btb_427 : _GEN_426; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_428 = 9'h1ac == io_ar_addr ? btb_428 : _GEN_427; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_429 = 9'h1ad == io_ar_addr ? btb_429 : _GEN_428; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_430 = 9'h1ae == io_ar_addr ? btb_430 : _GEN_429; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_431 = 9'h1af == io_ar_addr ? btb_431 : _GEN_430; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_432 = 9'h1b0 == io_ar_addr ? btb_432 : _GEN_431; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_433 = 9'h1b1 == io_ar_addr ? btb_433 : _GEN_432; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_434 = 9'h1b2 == io_ar_addr ? btb_434 : _GEN_433; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_435 = 9'h1b3 == io_ar_addr ? btb_435 : _GEN_434; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_436 = 9'h1b4 == io_ar_addr ? btb_436 : _GEN_435; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_437 = 9'h1b5 == io_ar_addr ? btb_437 : _GEN_436; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_438 = 9'h1b6 == io_ar_addr ? btb_438 : _GEN_437; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_439 = 9'h1b7 == io_ar_addr ? btb_439 : _GEN_438; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_440 = 9'h1b8 == io_ar_addr ? btb_440 : _GEN_439; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_441 = 9'h1b9 == io_ar_addr ? btb_441 : _GEN_440; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_442 = 9'h1ba == io_ar_addr ? btb_442 : _GEN_441; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_443 = 9'h1bb == io_ar_addr ? btb_443 : _GEN_442; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_444 = 9'h1bc == io_ar_addr ? btb_444 : _GEN_443; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_445 = 9'h1bd == io_ar_addr ? btb_445 : _GEN_444; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_446 = 9'h1be == io_ar_addr ? btb_446 : _GEN_445; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_447 = 9'h1bf == io_ar_addr ? btb_447 : _GEN_446; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_448 = 9'h1c0 == io_ar_addr ? btb_448 : _GEN_447; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_449 = 9'h1c1 == io_ar_addr ? btb_449 : _GEN_448; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_450 = 9'h1c2 == io_ar_addr ? btb_450 : _GEN_449; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_451 = 9'h1c3 == io_ar_addr ? btb_451 : _GEN_450; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_452 = 9'h1c4 == io_ar_addr ? btb_452 : _GEN_451; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_453 = 9'h1c5 == io_ar_addr ? btb_453 : _GEN_452; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_454 = 9'h1c6 == io_ar_addr ? btb_454 : _GEN_453; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_455 = 9'h1c7 == io_ar_addr ? btb_455 : _GEN_454; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_456 = 9'h1c8 == io_ar_addr ? btb_456 : _GEN_455; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_457 = 9'h1c9 == io_ar_addr ? btb_457 : _GEN_456; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_458 = 9'h1ca == io_ar_addr ? btb_458 : _GEN_457; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_459 = 9'h1cb == io_ar_addr ? btb_459 : _GEN_458; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_460 = 9'h1cc == io_ar_addr ? btb_460 : _GEN_459; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_461 = 9'h1cd == io_ar_addr ? btb_461 : _GEN_460; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_462 = 9'h1ce == io_ar_addr ? btb_462 : _GEN_461; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_463 = 9'h1cf == io_ar_addr ? btb_463 : _GEN_462; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_464 = 9'h1d0 == io_ar_addr ? btb_464 : _GEN_463; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_465 = 9'h1d1 == io_ar_addr ? btb_465 : _GEN_464; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_466 = 9'h1d2 == io_ar_addr ? btb_466 : _GEN_465; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_467 = 9'h1d3 == io_ar_addr ? btb_467 : _GEN_466; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_468 = 9'h1d4 == io_ar_addr ? btb_468 : _GEN_467; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_469 = 9'h1d5 == io_ar_addr ? btb_469 : _GEN_468; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_470 = 9'h1d6 == io_ar_addr ? btb_470 : _GEN_469; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_471 = 9'h1d7 == io_ar_addr ? btb_471 : _GEN_470; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_472 = 9'h1d8 == io_ar_addr ? btb_472 : _GEN_471; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_473 = 9'h1d9 == io_ar_addr ? btb_473 : _GEN_472; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_474 = 9'h1da == io_ar_addr ? btb_474 : _GEN_473; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_475 = 9'h1db == io_ar_addr ? btb_475 : _GEN_474; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_476 = 9'h1dc == io_ar_addr ? btb_476 : _GEN_475; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_477 = 9'h1dd == io_ar_addr ? btb_477 : _GEN_476; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_478 = 9'h1de == io_ar_addr ? btb_478 : _GEN_477; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_479 = 9'h1df == io_ar_addr ? btb_479 : _GEN_478; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_480 = 9'h1e0 == io_ar_addr ? btb_480 : _GEN_479; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_481 = 9'h1e1 == io_ar_addr ? btb_481 : _GEN_480; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_482 = 9'h1e2 == io_ar_addr ? btb_482 : _GEN_481; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_483 = 9'h1e3 == io_ar_addr ? btb_483 : _GEN_482; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_484 = 9'h1e4 == io_ar_addr ? btb_484 : _GEN_483; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_485 = 9'h1e5 == io_ar_addr ? btb_485 : _GEN_484; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_486 = 9'h1e6 == io_ar_addr ? btb_486 : _GEN_485; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_487 = 9'h1e7 == io_ar_addr ? btb_487 : _GEN_486; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_488 = 9'h1e8 == io_ar_addr ? btb_488 : _GEN_487; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_489 = 9'h1e9 == io_ar_addr ? btb_489 : _GEN_488; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_490 = 9'h1ea == io_ar_addr ? btb_490 : _GEN_489; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_491 = 9'h1eb == io_ar_addr ? btb_491 : _GEN_490; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_492 = 9'h1ec == io_ar_addr ? btb_492 : _GEN_491; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_493 = 9'h1ed == io_ar_addr ? btb_493 : _GEN_492; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_494 = 9'h1ee == io_ar_addr ? btb_494 : _GEN_493; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_495 = 9'h1ef == io_ar_addr ? btb_495 : _GEN_494; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_496 = 9'h1f0 == io_ar_addr ? btb_496 : _GEN_495; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_497 = 9'h1f1 == io_ar_addr ? btb_497 : _GEN_496; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_498 = 9'h1f2 == io_ar_addr ? btb_498 : _GEN_497; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_499 = 9'h1f3 == io_ar_addr ? btb_499 : _GEN_498; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_500 = 9'h1f4 == io_ar_addr ? btb_500 : _GEN_499; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_501 = 9'h1f5 == io_ar_addr ? btb_501 : _GEN_500; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_502 = 9'h1f6 == io_ar_addr ? btb_502 : _GEN_501; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_503 = 9'h1f7 == io_ar_addr ? btb_503 : _GEN_502; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_504 = 9'h1f8 == io_ar_addr ? btb_504 : _GEN_503; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_505 = 9'h1f9 == io_ar_addr ? btb_505 : _GEN_504; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_506 = 9'h1fa == io_ar_addr ? btb_506 : _GEN_505; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_507 = 9'h1fb == io_ar_addr ? btb_507 : _GEN_506; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_508 = 9'h1fc == io_ar_addr ? btb_508 : _GEN_507; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_509 = 9'h1fd == io_ar_addr ? btb_509 : _GEN_508; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_510 = 9'h1fe == io_ar_addr ? btb_510 : _GEN_509; // @[ports_lookup_table.scala 82:{12,12}]
  wire [7:0] _GEN_513 = 9'h1 == io_aw_addr ? btb_1 : btb_0; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_514 = 9'h2 == io_aw_addr ? btb_2 : _GEN_513; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_515 = 9'h3 == io_aw_addr ? btb_3 : _GEN_514; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_516 = 9'h4 == io_aw_addr ? btb_4 : _GEN_515; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_517 = 9'h5 == io_aw_addr ? btb_5 : _GEN_516; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_518 = 9'h6 == io_aw_addr ? btb_6 : _GEN_517; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_519 = 9'h7 == io_aw_addr ? btb_7 : _GEN_518; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_520 = 9'h8 == io_aw_addr ? btb_8 : _GEN_519; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_521 = 9'h9 == io_aw_addr ? btb_9 : _GEN_520; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_522 = 9'ha == io_aw_addr ? btb_10 : _GEN_521; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_523 = 9'hb == io_aw_addr ? btb_11 : _GEN_522; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_524 = 9'hc == io_aw_addr ? btb_12 : _GEN_523; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_525 = 9'hd == io_aw_addr ? btb_13 : _GEN_524; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_526 = 9'he == io_aw_addr ? btb_14 : _GEN_525; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_527 = 9'hf == io_aw_addr ? btb_15 : _GEN_526; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_528 = 9'h10 == io_aw_addr ? btb_16 : _GEN_527; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_529 = 9'h11 == io_aw_addr ? btb_17 : _GEN_528; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_530 = 9'h12 == io_aw_addr ? btb_18 : _GEN_529; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_531 = 9'h13 == io_aw_addr ? btb_19 : _GEN_530; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_532 = 9'h14 == io_aw_addr ? btb_20 : _GEN_531; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_533 = 9'h15 == io_aw_addr ? btb_21 : _GEN_532; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_534 = 9'h16 == io_aw_addr ? btb_22 : _GEN_533; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_535 = 9'h17 == io_aw_addr ? btb_23 : _GEN_534; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_536 = 9'h18 == io_aw_addr ? btb_24 : _GEN_535; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_537 = 9'h19 == io_aw_addr ? btb_25 : _GEN_536; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_538 = 9'h1a == io_aw_addr ? btb_26 : _GEN_537; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_539 = 9'h1b == io_aw_addr ? btb_27 : _GEN_538; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_540 = 9'h1c == io_aw_addr ? btb_28 : _GEN_539; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_541 = 9'h1d == io_aw_addr ? btb_29 : _GEN_540; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_542 = 9'h1e == io_aw_addr ? btb_30 : _GEN_541; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_543 = 9'h1f == io_aw_addr ? btb_31 : _GEN_542; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_544 = 9'h20 == io_aw_addr ? btb_32 : _GEN_543; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_545 = 9'h21 == io_aw_addr ? btb_33 : _GEN_544; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_546 = 9'h22 == io_aw_addr ? btb_34 : _GEN_545; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_547 = 9'h23 == io_aw_addr ? btb_35 : _GEN_546; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_548 = 9'h24 == io_aw_addr ? btb_36 : _GEN_547; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_549 = 9'h25 == io_aw_addr ? btb_37 : _GEN_548; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_550 = 9'h26 == io_aw_addr ? btb_38 : _GEN_549; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_551 = 9'h27 == io_aw_addr ? btb_39 : _GEN_550; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_552 = 9'h28 == io_aw_addr ? btb_40 : _GEN_551; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_553 = 9'h29 == io_aw_addr ? btb_41 : _GEN_552; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_554 = 9'h2a == io_aw_addr ? btb_42 : _GEN_553; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_555 = 9'h2b == io_aw_addr ? btb_43 : _GEN_554; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_556 = 9'h2c == io_aw_addr ? btb_44 : _GEN_555; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_557 = 9'h2d == io_aw_addr ? btb_45 : _GEN_556; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_558 = 9'h2e == io_aw_addr ? btb_46 : _GEN_557; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_559 = 9'h2f == io_aw_addr ? btb_47 : _GEN_558; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_560 = 9'h30 == io_aw_addr ? btb_48 : _GEN_559; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_561 = 9'h31 == io_aw_addr ? btb_49 : _GEN_560; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_562 = 9'h32 == io_aw_addr ? btb_50 : _GEN_561; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_563 = 9'h33 == io_aw_addr ? btb_51 : _GEN_562; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_564 = 9'h34 == io_aw_addr ? btb_52 : _GEN_563; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_565 = 9'h35 == io_aw_addr ? btb_53 : _GEN_564; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_566 = 9'h36 == io_aw_addr ? btb_54 : _GEN_565; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_567 = 9'h37 == io_aw_addr ? btb_55 : _GEN_566; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_568 = 9'h38 == io_aw_addr ? btb_56 : _GEN_567; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_569 = 9'h39 == io_aw_addr ? btb_57 : _GEN_568; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_570 = 9'h3a == io_aw_addr ? btb_58 : _GEN_569; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_571 = 9'h3b == io_aw_addr ? btb_59 : _GEN_570; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_572 = 9'h3c == io_aw_addr ? btb_60 : _GEN_571; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_573 = 9'h3d == io_aw_addr ? btb_61 : _GEN_572; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_574 = 9'h3e == io_aw_addr ? btb_62 : _GEN_573; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_575 = 9'h3f == io_aw_addr ? btb_63 : _GEN_574; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_576 = 9'h40 == io_aw_addr ? btb_64 : _GEN_575; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_577 = 9'h41 == io_aw_addr ? btb_65 : _GEN_576; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_578 = 9'h42 == io_aw_addr ? btb_66 : _GEN_577; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_579 = 9'h43 == io_aw_addr ? btb_67 : _GEN_578; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_580 = 9'h44 == io_aw_addr ? btb_68 : _GEN_579; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_581 = 9'h45 == io_aw_addr ? btb_69 : _GEN_580; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_582 = 9'h46 == io_aw_addr ? btb_70 : _GEN_581; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_583 = 9'h47 == io_aw_addr ? btb_71 : _GEN_582; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_584 = 9'h48 == io_aw_addr ? btb_72 : _GEN_583; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_585 = 9'h49 == io_aw_addr ? btb_73 : _GEN_584; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_586 = 9'h4a == io_aw_addr ? btb_74 : _GEN_585; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_587 = 9'h4b == io_aw_addr ? btb_75 : _GEN_586; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_588 = 9'h4c == io_aw_addr ? btb_76 : _GEN_587; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_589 = 9'h4d == io_aw_addr ? btb_77 : _GEN_588; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_590 = 9'h4e == io_aw_addr ? btb_78 : _GEN_589; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_591 = 9'h4f == io_aw_addr ? btb_79 : _GEN_590; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_592 = 9'h50 == io_aw_addr ? btb_80 : _GEN_591; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_593 = 9'h51 == io_aw_addr ? btb_81 : _GEN_592; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_594 = 9'h52 == io_aw_addr ? btb_82 : _GEN_593; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_595 = 9'h53 == io_aw_addr ? btb_83 : _GEN_594; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_596 = 9'h54 == io_aw_addr ? btb_84 : _GEN_595; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_597 = 9'h55 == io_aw_addr ? btb_85 : _GEN_596; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_598 = 9'h56 == io_aw_addr ? btb_86 : _GEN_597; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_599 = 9'h57 == io_aw_addr ? btb_87 : _GEN_598; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_600 = 9'h58 == io_aw_addr ? btb_88 : _GEN_599; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_601 = 9'h59 == io_aw_addr ? btb_89 : _GEN_600; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_602 = 9'h5a == io_aw_addr ? btb_90 : _GEN_601; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_603 = 9'h5b == io_aw_addr ? btb_91 : _GEN_602; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_604 = 9'h5c == io_aw_addr ? btb_92 : _GEN_603; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_605 = 9'h5d == io_aw_addr ? btb_93 : _GEN_604; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_606 = 9'h5e == io_aw_addr ? btb_94 : _GEN_605; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_607 = 9'h5f == io_aw_addr ? btb_95 : _GEN_606; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_608 = 9'h60 == io_aw_addr ? btb_96 : _GEN_607; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_609 = 9'h61 == io_aw_addr ? btb_97 : _GEN_608; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_610 = 9'h62 == io_aw_addr ? btb_98 : _GEN_609; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_611 = 9'h63 == io_aw_addr ? btb_99 : _GEN_610; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_612 = 9'h64 == io_aw_addr ? btb_100 : _GEN_611; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_613 = 9'h65 == io_aw_addr ? btb_101 : _GEN_612; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_614 = 9'h66 == io_aw_addr ? btb_102 : _GEN_613; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_615 = 9'h67 == io_aw_addr ? btb_103 : _GEN_614; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_616 = 9'h68 == io_aw_addr ? btb_104 : _GEN_615; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_617 = 9'h69 == io_aw_addr ? btb_105 : _GEN_616; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_618 = 9'h6a == io_aw_addr ? btb_106 : _GEN_617; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_619 = 9'h6b == io_aw_addr ? btb_107 : _GEN_618; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_620 = 9'h6c == io_aw_addr ? btb_108 : _GEN_619; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_621 = 9'h6d == io_aw_addr ? btb_109 : _GEN_620; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_622 = 9'h6e == io_aw_addr ? btb_110 : _GEN_621; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_623 = 9'h6f == io_aw_addr ? btb_111 : _GEN_622; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_624 = 9'h70 == io_aw_addr ? btb_112 : _GEN_623; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_625 = 9'h71 == io_aw_addr ? btb_113 : _GEN_624; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_626 = 9'h72 == io_aw_addr ? btb_114 : _GEN_625; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_627 = 9'h73 == io_aw_addr ? btb_115 : _GEN_626; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_628 = 9'h74 == io_aw_addr ? btb_116 : _GEN_627; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_629 = 9'h75 == io_aw_addr ? btb_117 : _GEN_628; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_630 = 9'h76 == io_aw_addr ? btb_118 : _GEN_629; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_631 = 9'h77 == io_aw_addr ? btb_119 : _GEN_630; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_632 = 9'h78 == io_aw_addr ? btb_120 : _GEN_631; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_633 = 9'h79 == io_aw_addr ? btb_121 : _GEN_632; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_634 = 9'h7a == io_aw_addr ? btb_122 : _GEN_633; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_635 = 9'h7b == io_aw_addr ? btb_123 : _GEN_634; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_636 = 9'h7c == io_aw_addr ? btb_124 : _GEN_635; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_637 = 9'h7d == io_aw_addr ? btb_125 : _GEN_636; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_638 = 9'h7e == io_aw_addr ? btb_126 : _GEN_637; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_639 = 9'h7f == io_aw_addr ? btb_127 : _GEN_638; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_640 = 9'h80 == io_aw_addr ? btb_128 : _GEN_639; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_641 = 9'h81 == io_aw_addr ? btb_129 : _GEN_640; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_642 = 9'h82 == io_aw_addr ? btb_130 : _GEN_641; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_643 = 9'h83 == io_aw_addr ? btb_131 : _GEN_642; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_644 = 9'h84 == io_aw_addr ? btb_132 : _GEN_643; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_645 = 9'h85 == io_aw_addr ? btb_133 : _GEN_644; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_646 = 9'h86 == io_aw_addr ? btb_134 : _GEN_645; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_647 = 9'h87 == io_aw_addr ? btb_135 : _GEN_646; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_648 = 9'h88 == io_aw_addr ? btb_136 : _GEN_647; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_649 = 9'h89 == io_aw_addr ? btb_137 : _GEN_648; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_650 = 9'h8a == io_aw_addr ? btb_138 : _GEN_649; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_651 = 9'h8b == io_aw_addr ? btb_139 : _GEN_650; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_652 = 9'h8c == io_aw_addr ? btb_140 : _GEN_651; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_653 = 9'h8d == io_aw_addr ? btb_141 : _GEN_652; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_654 = 9'h8e == io_aw_addr ? btb_142 : _GEN_653; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_655 = 9'h8f == io_aw_addr ? btb_143 : _GEN_654; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_656 = 9'h90 == io_aw_addr ? btb_144 : _GEN_655; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_657 = 9'h91 == io_aw_addr ? btb_145 : _GEN_656; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_658 = 9'h92 == io_aw_addr ? btb_146 : _GEN_657; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_659 = 9'h93 == io_aw_addr ? btb_147 : _GEN_658; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_660 = 9'h94 == io_aw_addr ? btb_148 : _GEN_659; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_661 = 9'h95 == io_aw_addr ? btb_149 : _GEN_660; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_662 = 9'h96 == io_aw_addr ? btb_150 : _GEN_661; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_663 = 9'h97 == io_aw_addr ? btb_151 : _GEN_662; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_664 = 9'h98 == io_aw_addr ? btb_152 : _GEN_663; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_665 = 9'h99 == io_aw_addr ? btb_153 : _GEN_664; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_666 = 9'h9a == io_aw_addr ? btb_154 : _GEN_665; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_667 = 9'h9b == io_aw_addr ? btb_155 : _GEN_666; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_668 = 9'h9c == io_aw_addr ? btb_156 : _GEN_667; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_669 = 9'h9d == io_aw_addr ? btb_157 : _GEN_668; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_670 = 9'h9e == io_aw_addr ? btb_158 : _GEN_669; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_671 = 9'h9f == io_aw_addr ? btb_159 : _GEN_670; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_672 = 9'ha0 == io_aw_addr ? btb_160 : _GEN_671; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_673 = 9'ha1 == io_aw_addr ? btb_161 : _GEN_672; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_674 = 9'ha2 == io_aw_addr ? btb_162 : _GEN_673; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_675 = 9'ha3 == io_aw_addr ? btb_163 : _GEN_674; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_676 = 9'ha4 == io_aw_addr ? btb_164 : _GEN_675; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_677 = 9'ha5 == io_aw_addr ? btb_165 : _GEN_676; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_678 = 9'ha6 == io_aw_addr ? btb_166 : _GEN_677; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_679 = 9'ha7 == io_aw_addr ? btb_167 : _GEN_678; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_680 = 9'ha8 == io_aw_addr ? btb_168 : _GEN_679; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_681 = 9'ha9 == io_aw_addr ? btb_169 : _GEN_680; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_682 = 9'haa == io_aw_addr ? btb_170 : _GEN_681; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_683 = 9'hab == io_aw_addr ? btb_171 : _GEN_682; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_684 = 9'hac == io_aw_addr ? btb_172 : _GEN_683; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_685 = 9'had == io_aw_addr ? btb_173 : _GEN_684; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_686 = 9'hae == io_aw_addr ? btb_174 : _GEN_685; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_687 = 9'haf == io_aw_addr ? btb_175 : _GEN_686; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_688 = 9'hb0 == io_aw_addr ? btb_176 : _GEN_687; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_689 = 9'hb1 == io_aw_addr ? btb_177 : _GEN_688; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_690 = 9'hb2 == io_aw_addr ? btb_178 : _GEN_689; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_691 = 9'hb3 == io_aw_addr ? btb_179 : _GEN_690; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_692 = 9'hb4 == io_aw_addr ? btb_180 : _GEN_691; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_693 = 9'hb5 == io_aw_addr ? btb_181 : _GEN_692; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_694 = 9'hb6 == io_aw_addr ? btb_182 : _GEN_693; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_695 = 9'hb7 == io_aw_addr ? btb_183 : _GEN_694; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_696 = 9'hb8 == io_aw_addr ? btb_184 : _GEN_695; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_697 = 9'hb9 == io_aw_addr ? btb_185 : _GEN_696; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_698 = 9'hba == io_aw_addr ? btb_186 : _GEN_697; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_699 = 9'hbb == io_aw_addr ? btb_187 : _GEN_698; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_700 = 9'hbc == io_aw_addr ? btb_188 : _GEN_699; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_701 = 9'hbd == io_aw_addr ? btb_189 : _GEN_700; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_702 = 9'hbe == io_aw_addr ? btb_190 : _GEN_701; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_703 = 9'hbf == io_aw_addr ? btb_191 : _GEN_702; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_704 = 9'hc0 == io_aw_addr ? btb_192 : _GEN_703; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_705 = 9'hc1 == io_aw_addr ? btb_193 : _GEN_704; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_706 = 9'hc2 == io_aw_addr ? btb_194 : _GEN_705; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_707 = 9'hc3 == io_aw_addr ? btb_195 : _GEN_706; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_708 = 9'hc4 == io_aw_addr ? btb_196 : _GEN_707; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_709 = 9'hc5 == io_aw_addr ? btb_197 : _GEN_708; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_710 = 9'hc6 == io_aw_addr ? btb_198 : _GEN_709; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_711 = 9'hc7 == io_aw_addr ? btb_199 : _GEN_710; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_712 = 9'hc8 == io_aw_addr ? btb_200 : _GEN_711; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_713 = 9'hc9 == io_aw_addr ? btb_201 : _GEN_712; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_714 = 9'hca == io_aw_addr ? btb_202 : _GEN_713; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_715 = 9'hcb == io_aw_addr ? btb_203 : _GEN_714; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_716 = 9'hcc == io_aw_addr ? btb_204 : _GEN_715; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_717 = 9'hcd == io_aw_addr ? btb_205 : _GEN_716; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_718 = 9'hce == io_aw_addr ? btb_206 : _GEN_717; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_719 = 9'hcf == io_aw_addr ? btb_207 : _GEN_718; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_720 = 9'hd0 == io_aw_addr ? btb_208 : _GEN_719; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_721 = 9'hd1 == io_aw_addr ? btb_209 : _GEN_720; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_722 = 9'hd2 == io_aw_addr ? btb_210 : _GEN_721; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_723 = 9'hd3 == io_aw_addr ? btb_211 : _GEN_722; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_724 = 9'hd4 == io_aw_addr ? btb_212 : _GEN_723; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_725 = 9'hd5 == io_aw_addr ? btb_213 : _GEN_724; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_726 = 9'hd6 == io_aw_addr ? btb_214 : _GEN_725; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_727 = 9'hd7 == io_aw_addr ? btb_215 : _GEN_726; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_728 = 9'hd8 == io_aw_addr ? btb_216 : _GEN_727; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_729 = 9'hd9 == io_aw_addr ? btb_217 : _GEN_728; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_730 = 9'hda == io_aw_addr ? btb_218 : _GEN_729; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_731 = 9'hdb == io_aw_addr ? btb_219 : _GEN_730; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_732 = 9'hdc == io_aw_addr ? btb_220 : _GEN_731; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_733 = 9'hdd == io_aw_addr ? btb_221 : _GEN_732; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_734 = 9'hde == io_aw_addr ? btb_222 : _GEN_733; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_735 = 9'hdf == io_aw_addr ? btb_223 : _GEN_734; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_736 = 9'he0 == io_aw_addr ? btb_224 : _GEN_735; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_737 = 9'he1 == io_aw_addr ? btb_225 : _GEN_736; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_738 = 9'he2 == io_aw_addr ? btb_226 : _GEN_737; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_739 = 9'he3 == io_aw_addr ? btb_227 : _GEN_738; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_740 = 9'he4 == io_aw_addr ? btb_228 : _GEN_739; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_741 = 9'he5 == io_aw_addr ? btb_229 : _GEN_740; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_742 = 9'he6 == io_aw_addr ? btb_230 : _GEN_741; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_743 = 9'he7 == io_aw_addr ? btb_231 : _GEN_742; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_744 = 9'he8 == io_aw_addr ? btb_232 : _GEN_743; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_745 = 9'he9 == io_aw_addr ? btb_233 : _GEN_744; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_746 = 9'hea == io_aw_addr ? btb_234 : _GEN_745; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_747 = 9'heb == io_aw_addr ? btb_235 : _GEN_746; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_748 = 9'hec == io_aw_addr ? btb_236 : _GEN_747; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_749 = 9'hed == io_aw_addr ? btb_237 : _GEN_748; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_750 = 9'hee == io_aw_addr ? btb_238 : _GEN_749; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_751 = 9'hef == io_aw_addr ? btb_239 : _GEN_750; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_752 = 9'hf0 == io_aw_addr ? btb_240 : _GEN_751; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_753 = 9'hf1 == io_aw_addr ? btb_241 : _GEN_752; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_754 = 9'hf2 == io_aw_addr ? btb_242 : _GEN_753; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_755 = 9'hf3 == io_aw_addr ? btb_243 : _GEN_754; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_756 = 9'hf4 == io_aw_addr ? btb_244 : _GEN_755; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_757 = 9'hf5 == io_aw_addr ? btb_245 : _GEN_756; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_758 = 9'hf6 == io_aw_addr ? btb_246 : _GEN_757; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_759 = 9'hf7 == io_aw_addr ? btb_247 : _GEN_758; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_760 = 9'hf8 == io_aw_addr ? btb_248 : _GEN_759; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_761 = 9'hf9 == io_aw_addr ? btb_249 : _GEN_760; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_762 = 9'hfa == io_aw_addr ? btb_250 : _GEN_761; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_763 = 9'hfb == io_aw_addr ? btb_251 : _GEN_762; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_764 = 9'hfc == io_aw_addr ? btb_252 : _GEN_763; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_765 = 9'hfd == io_aw_addr ? btb_253 : _GEN_764; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_766 = 9'hfe == io_aw_addr ? btb_254 : _GEN_765; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_767 = 9'hff == io_aw_addr ? btb_255 : _GEN_766; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_768 = 9'h100 == io_aw_addr ? btb_256 : _GEN_767; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_769 = 9'h101 == io_aw_addr ? btb_257 : _GEN_768; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_770 = 9'h102 == io_aw_addr ? btb_258 : _GEN_769; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_771 = 9'h103 == io_aw_addr ? btb_259 : _GEN_770; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_772 = 9'h104 == io_aw_addr ? btb_260 : _GEN_771; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_773 = 9'h105 == io_aw_addr ? btb_261 : _GEN_772; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_774 = 9'h106 == io_aw_addr ? btb_262 : _GEN_773; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_775 = 9'h107 == io_aw_addr ? btb_263 : _GEN_774; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_776 = 9'h108 == io_aw_addr ? btb_264 : _GEN_775; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_777 = 9'h109 == io_aw_addr ? btb_265 : _GEN_776; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_778 = 9'h10a == io_aw_addr ? btb_266 : _GEN_777; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_779 = 9'h10b == io_aw_addr ? btb_267 : _GEN_778; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_780 = 9'h10c == io_aw_addr ? btb_268 : _GEN_779; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_781 = 9'h10d == io_aw_addr ? btb_269 : _GEN_780; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_782 = 9'h10e == io_aw_addr ? btb_270 : _GEN_781; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_783 = 9'h10f == io_aw_addr ? btb_271 : _GEN_782; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_784 = 9'h110 == io_aw_addr ? btb_272 : _GEN_783; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_785 = 9'h111 == io_aw_addr ? btb_273 : _GEN_784; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_786 = 9'h112 == io_aw_addr ? btb_274 : _GEN_785; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_787 = 9'h113 == io_aw_addr ? btb_275 : _GEN_786; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_788 = 9'h114 == io_aw_addr ? btb_276 : _GEN_787; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_789 = 9'h115 == io_aw_addr ? btb_277 : _GEN_788; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_790 = 9'h116 == io_aw_addr ? btb_278 : _GEN_789; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_791 = 9'h117 == io_aw_addr ? btb_279 : _GEN_790; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_792 = 9'h118 == io_aw_addr ? btb_280 : _GEN_791; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_793 = 9'h119 == io_aw_addr ? btb_281 : _GEN_792; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_794 = 9'h11a == io_aw_addr ? btb_282 : _GEN_793; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_795 = 9'h11b == io_aw_addr ? btb_283 : _GEN_794; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_796 = 9'h11c == io_aw_addr ? btb_284 : _GEN_795; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_797 = 9'h11d == io_aw_addr ? btb_285 : _GEN_796; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_798 = 9'h11e == io_aw_addr ? btb_286 : _GEN_797; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_799 = 9'h11f == io_aw_addr ? btb_287 : _GEN_798; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_800 = 9'h120 == io_aw_addr ? btb_288 : _GEN_799; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_801 = 9'h121 == io_aw_addr ? btb_289 : _GEN_800; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_802 = 9'h122 == io_aw_addr ? btb_290 : _GEN_801; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_803 = 9'h123 == io_aw_addr ? btb_291 : _GEN_802; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_804 = 9'h124 == io_aw_addr ? btb_292 : _GEN_803; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_805 = 9'h125 == io_aw_addr ? btb_293 : _GEN_804; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_806 = 9'h126 == io_aw_addr ? btb_294 : _GEN_805; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_807 = 9'h127 == io_aw_addr ? btb_295 : _GEN_806; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_808 = 9'h128 == io_aw_addr ? btb_296 : _GEN_807; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_809 = 9'h129 == io_aw_addr ? btb_297 : _GEN_808; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_810 = 9'h12a == io_aw_addr ? btb_298 : _GEN_809; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_811 = 9'h12b == io_aw_addr ? btb_299 : _GEN_810; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_812 = 9'h12c == io_aw_addr ? btb_300 : _GEN_811; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_813 = 9'h12d == io_aw_addr ? btb_301 : _GEN_812; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_814 = 9'h12e == io_aw_addr ? btb_302 : _GEN_813; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_815 = 9'h12f == io_aw_addr ? btb_303 : _GEN_814; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_816 = 9'h130 == io_aw_addr ? btb_304 : _GEN_815; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_817 = 9'h131 == io_aw_addr ? btb_305 : _GEN_816; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_818 = 9'h132 == io_aw_addr ? btb_306 : _GEN_817; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_819 = 9'h133 == io_aw_addr ? btb_307 : _GEN_818; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_820 = 9'h134 == io_aw_addr ? btb_308 : _GEN_819; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_821 = 9'h135 == io_aw_addr ? btb_309 : _GEN_820; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_822 = 9'h136 == io_aw_addr ? btb_310 : _GEN_821; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_823 = 9'h137 == io_aw_addr ? btb_311 : _GEN_822; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_824 = 9'h138 == io_aw_addr ? btb_312 : _GEN_823; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_825 = 9'h139 == io_aw_addr ? btb_313 : _GEN_824; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_826 = 9'h13a == io_aw_addr ? btb_314 : _GEN_825; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_827 = 9'h13b == io_aw_addr ? btb_315 : _GEN_826; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_828 = 9'h13c == io_aw_addr ? btb_316 : _GEN_827; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_829 = 9'h13d == io_aw_addr ? btb_317 : _GEN_828; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_830 = 9'h13e == io_aw_addr ? btb_318 : _GEN_829; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_831 = 9'h13f == io_aw_addr ? btb_319 : _GEN_830; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_832 = 9'h140 == io_aw_addr ? btb_320 : _GEN_831; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_833 = 9'h141 == io_aw_addr ? btb_321 : _GEN_832; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_834 = 9'h142 == io_aw_addr ? btb_322 : _GEN_833; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_835 = 9'h143 == io_aw_addr ? btb_323 : _GEN_834; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_836 = 9'h144 == io_aw_addr ? btb_324 : _GEN_835; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_837 = 9'h145 == io_aw_addr ? btb_325 : _GEN_836; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_838 = 9'h146 == io_aw_addr ? btb_326 : _GEN_837; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_839 = 9'h147 == io_aw_addr ? btb_327 : _GEN_838; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_840 = 9'h148 == io_aw_addr ? btb_328 : _GEN_839; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_841 = 9'h149 == io_aw_addr ? btb_329 : _GEN_840; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_842 = 9'h14a == io_aw_addr ? btb_330 : _GEN_841; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_843 = 9'h14b == io_aw_addr ? btb_331 : _GEN_842; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_844 = 9'h14c == io_aw_addr ? btb_332 : _GEN_843; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_845 = 9'h14d == io_aw_addr ? btb_333 : _GEN_844; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_846 = 9'h14e == io_aw_addr ? btb_334 : _GEN_845; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_847 = 9'h14f == io_aw_addr ? btb_335 : _GEN_846; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_848 = 9'h150 == io_aw_addr ? btb_336 : _GEN_847; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_849 = 9'h151 == io_aw_addr ? btb_337 : _GEN_848; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_850 = 9'h152 == io_aw_addr ? btb_338 : _GEN_849; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_851 = 9'h153 == io_aw_addr ? btb_339 : _GEN_850; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_852 = 9'h154 == io_aw_addr ? btb_340 : _GEN_851; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_853 = 9'h155 == io_aw_addr ? btb_341 : _GEN_852; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_854 = 9'h156 == io_aw_addr ? btb_342 : _GEN_853; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_855 = 9'h157 == io_aw_addr ? btb_343 : _GEN_854; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_856 = 9'h158 == io_aw_addr ? btb_344 : _GEN_855; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_857 = 9'h159 == io_aw_addr ? btb_345 : _GEN_856; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_858 = 9'h15a == io_aw_addr ? btb_346 : _GEN_857; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_859 = 9'h15b == io_aw_addr ? btb_347 : _GEN_858; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_860 = 9'h15c == io_aw_addr ? btb_348 : _GEN_859; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_861 = 9'h15d == io_aw_addr ? btb_349 : _GEN_860; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_862 = 9'h15e == io_aw_addr ? btb_350 : _GEN_861; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_863 = 9'h15f == io_aw_addr ? btb_351 : _GEN_862; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_864 = 9'h160 == io_aw_addr ? btb_352 : _GEN_863; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_865 = 9'h161 == io_aw_addr ? btb_353 : _GEN_864; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_866 = 9'h162 == io_aw_addr ? btb_354 : _GEN_865; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_867 = 9'h163 == io_aw_addr ? btb_355 : _GEN_866; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_868 = 9'h164 == io_aw_addr ? btb_356 : _GEN_867; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_869 = 9'h165 == io_aw_addr ? btb_357 : _GEN_868; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_870 = 9'h166 == io_aw_addr ? btb_358 : _GEN_869; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_871 = 9'h167 == io_aw_addr ? btb_359 : _GEN_870; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_872 = 9'h168 == io_aw_addr ? btb_360 : _GEN_871; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_873 = 9'h169 == io_aw_addr ? btb_361 : _GEN_872; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_874 = 9'h16a == io_aw_addr ? btb_362 : _GEN_873; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_875 = 9'h16b == io_aw_addr ? btb_363 : _GEN_874; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_876 = 9'h16c == io_aw_addr ? btb_364 : _GEN_875; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_877 = 9'h16d == io_aw_addr ? btb_365 : _GEN_876; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_878 = 9'h16e == io_aw_addr ? btb_366 : _GEN_877; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_879 = 9'h16f == io_aw_addr ? btb_367 : _GEN_878; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_880 = 9'h170 == io_aw_addr ? btb_368 : _GEN_879; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_881 = 9'h171 == io_aw_addr ? btb_369 : _GEN_880; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_882 = 9'h172 == io_aw_addr ? btb_370 : _GEN_881; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_883 = 9'h173 == io_aw_addr ? btb_371 : _GEN_882; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_884 = 9'h174 == io_aw_addr ? btb_372 : _GEN_883; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_885 = 9'h175 == io_aw_addr ? btb_373 : _GEN_884; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_886 = 9'h176 == io_aw_addr ? btb_374 : _GEN_885; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_887 = 9'h177 == io_aw_addr ? btb_375 : _GEN_886; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_888 = 9'h178 == io_aw_addr ? btb_376 : _GEN_887; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_889 = 9'h179 == io_aw_addr ? btb_377 : _GEN_888; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_890 = 9'h17a == io_aw_addr ? btb_378 : _GEN_889; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_891 = 9'h17b == io_aw_addr ? btb_379 : _GEN_890; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_892 = 9'h17c == io_aw_addr ? btb_380 : _GEN_891; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_893 = 9'h17d == io_aw_addr ? btb_381 : _GEN_892; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_894 = 9'h17e == io_aw_addr ? btb_382 : _GEN_893; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_895 = 9'h17f == io_aw_addr ? btb_383 : _GEN_894; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_896 = 9'h180 == io_aw_addr ? btb_384 : _GEN_895; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_897 = 9'h181 == io_aw_addr ? btb_385 : _GEN_896; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_898 = 9'h182 == io_aw_addr ? btb_386 : _GEN_897; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_899 = 9'h183 == io_aw_addr ? btb_387 : _GEN_898; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_900 = 9'h184 == io_aw_addr ? btb_388 : _GEN_899; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_901 = 9'h185 == io_aw_addr ? btb_389 : _GEN_900; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_902 = 9'h186 == io_aw_addr ? btb_390 : _GEN_901; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_903 = 9'h187 == io_aw_addr ? btb_391 : _GEN_902; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_904 = 9'h188 == io_aw_addr ? btb_392 : _GEN_903; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_905 = 9'h189 == io_aw_addr ? btb_393 : _GEN_904; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_906 = 9'h18a == io_aw_addr ? btb_394 : _GEN_905; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_907 = 9'h18b == io_aw_addr ? btb_395 : _GEN_906; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_908 = 9'h18c == io_aw_addr ? btb_396 : _GEN_907; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_909 = 9'h18d == io_aw_addr ? btb_397 : _GEN_908; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_910 = 9'h18e == io_aw_addr ? btb_398 : _GEN_909; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_911 = 9'h18f == io_aw_addr ? btb_399 : _GEN_910; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_912 = 9'h190 == io_aw_addr ? btb_400 : _GEN_911; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_913 = 9'h191 == io_aw_addr ? btb_401 : _GEN_912; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_914 = 9'h192 == io_aw_addr ? btb_402 : _GEN_913; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_915 = 9'h193 == io_aw_addr ? btb_403 : _GEN_914; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_916 = 9'h194 == io_aw_addr ? btb_404 : _GEN_915; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_917 = 9'h195 == io_aw_addr ? btb_405 : _GEN_916; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_918 = 9'h196 == io_aw_addr ? btb_406 : _GEN_917; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_919 = 9'h197 == io_aw_addr ? btb_407 : _GEN_918; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_920 = 9'h198 == io_aw_addr ? btb_408 : _GEN_919; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_921 = 9'h199 == io_aw_addr ? btb_409 : _GEN_920; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_922 = 9'h19a == io_aw_addr ? btb_410 : _GEN_921; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_923 = 9'h19b == io_aw_addr ? btb_411 : _GEN_922; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_924 = 9'h19c == io_aw_addr ? btb_412 : _GEN_923; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_925 = 9'h19d == io_aw_addr ? btb_413 : _GEN_924; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_926 = 9'h19e == io_aw_addr ? btb_414 : _GEN_925; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_927 = 9'h19f == io_aw_addr ? btb_415 : _GEN_926; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_928 = 9'h1a0 == io_aw_addr ? btb_416 : _GEN_927; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_929 = 9'h1a1 == io_aw_addr ? btb_417 : _GEN_928; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_930 = 9'h1a2 == io_aw_addr ? btb_418 : _GEN_929; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_931 = 9'h1a3 == io_aw_addr ? btb_419 : _GEN_930; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_932 = 9'h1a4 == io_aw_addr ? btb_420 : _GEN_931; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_933 = 9'h1a5 == io_aw_addr ? btb_421 : _GEN_932; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_934 = 9'h1a6 == io_aw_addr ? btb_422 : _GEN_933; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_935 = 9'h1a7 == io_aw_addr ? btb_423 : _GEN_934; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_936 = 9'h1a8 == io_aw_addr ? btb_424 : _GEN_935; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_937 = 9'h1a9 == io_aw_addr ? btb_425 : _GEN_936; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_938 = 9'h1aa == io_aw_addr ? btb_426 : _GEN_937; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_939 = 9'h1ab == io_aw_addr ? btb_427 : _GEN_938; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_940 = 9'h1ac == io_aw_addr ? btb_428 : _GEN_939; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_941 = 9'h1ad == io_aw_addr ? btb_429 : _GEN_940; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_942 = 9'h1ae == io_aw_addr ? btb_430 : _GEN_941; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_943 = 9'h1af == io_aw_addr ? btb_431 : _GEN_942; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_944 = 9'h1b0 == io_aw_addr ? btb_432 : _GEN_943; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_945 = 9'h1b1 == io_aw_addr ? btb_433 : _GEN_944; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_946 = 9'h1b2 == io_aw_addr ? btb_434 : _GEN_945; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_947 = 9'h1b3 == io_aw_addr ? btb_435 : _GEN_946; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_948 = 9'h1b4 == io_aw_addr ? btb_436 : _GEN_947; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_949 = 9'h1b5 == io_aw_addr ? btb_437 : _GEN_948; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_950 = 9'h1b6 == io_aw_addr ? btb_438 : _GEN_949; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_951 = 9'h1b7 == io_aw_addr ? btb_439 : _GEN_950; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_952 = 9'h1b8 == io_aw_addr ? btb_440 : _GEN_951; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_953 = 9'h1b9 == io_aw_addr ? btb_441 : _GEN_952; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_954 = 9'h1ba == io_aw_addr ? btb_442 : _GEN_953; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_955 = 9'h1bb == io_aw_addr ? btb_443 : _GEN_954; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_956 = 9'h1bc == io_aw_addr ? btb_444 : _GEN_955; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_957 = 9'h1bd == io_aw_addr ? btb_445 : _GEN_956; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_958 = 9'h1be == io_aw_addr ? btb_446 : _GEN_957; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_959 = 9'h1bf == io_aw_addr ? btb_447 : _GEN_958; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_960 = 9'h1c0 == io_aw_addr ? btb_448 : _GEN_959; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_961 = 9'h1c1 == io_aw_addr ? btb_449 : _GEN_960; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_962 = 9'h1c2 == io_aw_addr ? btb_450 : _GEN_961; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_963 = 9'h1c3 == io_aw_addr ? btb_451 : _GEN_962; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_964 = 9'h1c4 == io_aw_addr ? btb_452 : _GEN_963; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_965 = 9'h1c5 == io_aw_addr ? btb_453 : _GEN_964; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_966 = 9'h1c6 == io_aw_addr ? btb_454 : _GEN_965; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_967 = 9'h1c7 == io_aw_addr ? btb_455 : _GEN_966; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_968 = 9'h1c8 == io_aw_addr ? btb_456 : _GEN_967; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_969 = 9'h1c9 == io_aw_addr ? btb_457 : _GEN_968; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_970 = 9'h1ca == io_aw_addr ? btb_458 : _GEN_969; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_971 = 9'h1cb == io_aw_addr ? btb_459 : _GEN_970; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_972 = 9'h1cc == io_aw_addr ? btb_460 : _GEN_971; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_973 = 9'h1cd == io_aw_addr ? btb_461 : _GEN_972; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_974 = 9'h1ce == io_aw_addr ? btb_462 : _GEN_973; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_975 = 9'h1cf == io_aw_addr ? btb_463 : _GEN_974; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_976 = 9'h1d0 == io_aw_addr ? btb_464 : _GEN_975; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_977 = 9'h1d1 == io_aw_addr ? btb_465 : _GEN_976; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_978 = 9'h1d2 == io_aw_addr ? btb_466 : _GEN_977; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_979 = 9'h1d3 == io_aw_addr ? btb_467 : _GEN_978; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_980 = 9'h1d4 == io_aw_addr ? btb_468 : _GEN_979; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_981 = 9'h1d5 == io_aw_addr ? btb_469 : _GEN_980; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_982 = 9'h1d6 == io_aw_addr ? btb_470 : _GEN_981; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_983 = 9'h1d7 == io_aw_addr ? btb_471 : _GEN_982; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_984 = 9'h1d8 == io_aw_addr ? btb_472 : _GEN_983; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_985 = 9'h1d9 == io_aw_addr ? btb_473 : _GEN_984; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_986 = 9'h1da == io_aw_addr ? btb_474 : _GEN_985; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_987 = 9'h1db == io_aw_addr ? btb_475 : _GEN_986; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_988 = 9'h1dc == io_aw_addr ? btb_476 : _GEN_987; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_989 = 9'h1dd == io_aw_addr ? btb_477 : _GEN_988; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_990 = 9'h1de == io_aw_addr ? btb_478 : _GEN_989; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_991 = 9'h1df == io_aw_addr ? btb_479 : _GEN_990; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_992 = 9'h1e0 == io_aw_addr ? btb_480 : _GEN_991; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_993 = 9'h1e1 == io_aw_addr ? btb_481 : _GEN_992; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_994 = 9'h1e2 == io_aw_addr ? btb_482 : _GEN_993; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_995 = 9'h1e3 == io_aw_addr ? btb_483 : _GEN_994; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_996 = 9'h1e4 == io_aw_addr ? btb_484 : _GEN_995; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_997 = 9'h1e5 == io_aw_addr ? btb_485 : _GEN_996; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_998 = 9'h1e6 == io_aw_addr ? btb_486 : _GEN_997; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_999 = 9'h1e7 == io_aw_addr ? btb_487 : _GEN_998; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1000 = 9'h1e8 == io_aw_addr ? btb_488 : _GEN_999; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1001 = 9'h1e9 == io_aw_addr ? btb_489 : _GEN_1000; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1002 = 9'h1ea == io_aw_addr ? btb_490 : _GEN_1001; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1003 = 9'h1eb == io_aw_addr ? btb_491 : _GEN_1002; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1004 = 9'h1ec == io_aw_addr ? btb_492 : _GEN_1003; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1005 = 9'h1ed == io_aw_addr ? btb_493 : _GEN_1004; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1006 = 9'h1ee == io_aw_addr ? btb_494 : _GEN_1005; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1007 = 9'h1ef == io_aw_addr ? btb_495 : _GEN_1006; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1008 = 9'h1f0 == io_aw_addr ? btb_496 : _GEN_1007; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1009 = 9'h1f1 == io_aw_addr ? btb_497 : _GEN_1008; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1010 = 9'h1f2 == io_aw_addr ? btb_498 : _GEN_1009; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1011 = 9'h1f3 == io_aw_addr ? btb_499 : _GEN_1010; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1012 = 9'h1f4 == io_aw_addr ? btb_500 : _GEN_1011; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1013 = 9'h1f5 == io_aw_addr ? btb_501 : _GEN_1012; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1014 = 9'h1f6 == io_aw_addr ? btb_502 : _GEN_1013; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1015 = 9'h1f7 == io_aw_addr ? btb_503 : _GEN_1014; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1016 = 9'h1f8 == io_aw_addr ? btb_504 : _GEN_1015; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1017 = 9'h1f9 == io_aw_addr ? btb_505 : _GEN_1016; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1018 = 9'h1fa == io_aw_addr ? btb_506 : _GEN_1017; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1019 = 9'h1fb == io_aw_addr ? btb_507 : _GEN_1018; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1020 = 9'h1fc == io_aw_addr ? btb_508 : _GEN_1019; // @[ports_lookup_table.scala 83:{27,27}]
  wire [7:0] _GEN_1021 = 9'h1fd == io_aw_addr ? btb_509 : _GEN_1020; // @[ports_lookup_table.scala 83:{27,27}]
  assign io_out = 9'h1ff == io_ar_addr ? btb_511 : _GEN_510; // @[ports_lookup_table.scala 82:{12,12}]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_0 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_0 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_0 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_0 <= btb_510;
      end else begin
        btb_0 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_1 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_1 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_1 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_1 <= btb_510;
      end else begin
        btb_1 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_2 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_2 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_2 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_2 <= btb_510;
      end else begin
        btb_2 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_3 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_3 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_3 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_3 <= btb_510;
      end else begin
        btb_3 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_4 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_4 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_4 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_4 <= btb_510;
      end else begin
        btb_4 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_5 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_5 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_5 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_5 <= btb_510;
      end else begin
        btb_5 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_6 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_6 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_6 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_6 <= btb_510;
      end else begin
        btb_6 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_7 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_7 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_7 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_7 <= btb_510;
      end else begin
        btb_7 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_8 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_8 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_8 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_8 <= btb_510;
      end else begin
        btb_8 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_9 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_9 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_9 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_9 <= btb_510;
      end else begin
        btb_9 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_10 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_10 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_10 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_10 <= btb_510;
      end else begin
        btb_10 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_11 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_11 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_11 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_11 <= btb_510;
      end else begin
        btb_11 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_12 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_12 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_12 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_12 <= btb_510;
      end else begin
        btb_12 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_13 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_13 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_13 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_13 <= btb_510;
      end else begin
        btb_13 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_14 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_14 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_14 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_14 <= btb_510;
      end else begin
        btb_14 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_15 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_15 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_15 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_15 <= btb_510;
      end else begin
        btb_15 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_16 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h10 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_16 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_16 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_16 <= btb_510;
      end else begin
        btb_16 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_17 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h11 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_17 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_17 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_17 <= btb_510;
      end else begin
        btb_17 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_18 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h12 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_18 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_18 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_18 <= btb_510;
      end else begin
        btb_18 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_19 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h13 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_19 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_19 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_19 <= btb_510;
      end else begin
        btb_19 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_20 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h14 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_20 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_20 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_20 <= btb_510;
      end else begin
        btb_20 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_21 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h15 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_21 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_21 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_21 <= btb_510;
      end else begin
        btb_21 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_22 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h16 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_22 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_22 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_22 <= btb_510;
      end else begin
        btb_22 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_23 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h17 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_23 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_23 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_23 <= btb_510;
      end else begin
        btb_23 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_24 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h18 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_24 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_24 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_24 <= btb_510;
      end else begin
        btb_24 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_25 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h19 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_25 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_25 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_25 <= btb_510;
      end else begin
        btb_25 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_26 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_26 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_26 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_26 <= btb_510;
      end else begin
        btb_26 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_27 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_27 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_27 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_27 <= btb_510;
      end else begin
        btb_27 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_28 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_28 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_28 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_28 <= btb_510;
      end else begin
        btb_28 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_29 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_29 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_29 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_29 <= btb_510;
      end else begin
        btb_29 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_30 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_30 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_30 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_30 <= btb_510;
      end else begin
        btb_30 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_31 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_31 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_31 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_31 <= btb_510;
      end else begin
        btb_31 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_32 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h20 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_32 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_32 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_32 <= btb_510;
      end else begin
        btb_32 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_33 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h21 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_33 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_33 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_33 <= btb_510;
      end else begin
        btb_33 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_34 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h22 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_34 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_34 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_34 <= btb_510;
      end else begin
        btb_34 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_35 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h23 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_35 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_35 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_35 <= btb_510;
      end else begin
        btb_35 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_36 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h24 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_36 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_36 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_36 <= btb_510;
      end else begin
        btb_36 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_37 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h25 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_37 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_37 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_37 <= btb_510;
      end else begin
        btb_37 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_38 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h26 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_38 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_38 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_38 <= btb_510;
      end else begin
        btb_38 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_39 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h27 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_39 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_39 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_39 <= btb_510;
      end else begin
        btb_39 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_40 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h28 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_40 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_40 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_40 <= btb_510;
      end else begin
        btb_40 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_41 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h29 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_41 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_41 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_41 <= btb_510;
      end else begin
        btb_41 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_42 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h2a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_42 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_42 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_42 <= btb_510;
      end else begin
        btb_42 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_43 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h2b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_43 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_43 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_43 <= btb_510;
      end else begin
        btb_43 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_44 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h2c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_44 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_44 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_44 <= btb_510;
      end else begin
        btb_44 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_45 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h2d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_45 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_45 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_45 <= btb_510;
      end else begin
        btb_45 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_46 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h2e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_46 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_46 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_46 <= btb_510;
      end else begin
        btb_46 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_47 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h2f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_47 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_47 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_47 <= btb_510;
      end else begin
        btb_47 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_48 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h30 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_48 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_48 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_48 <= btb_510;
      end else begin
        btb_48 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_49 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h31 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_49 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_49 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_49 <= btb_510;
      end else begin
        btb_49 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_50 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h32 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_50 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_50 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_50 <= btb_510;
      end else begin
        btb_50 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_51 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h33 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_51 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_51 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_51 <= btb_510;
      end else begin
        btb_51 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_52 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h34 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_52 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_52 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_52 <= btb_510;
      end else begin
        btb_52 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_53 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h35 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_53 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_53 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_53 <= btb_510;
      end else begin
        btb_53 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_54 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h36 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_54 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_54 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_54 <= btb_510;
      end else begin
        btb_54 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_55 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h37 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_55 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_55 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_55 <= btb_510;
      end else begin
        btb_55 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_56 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h38 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_56 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_56 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_56 <= btb_510;
      end else begin
        btb_56 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_57 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h39 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_57 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_57 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_57 <= btb_510;
      end else begin
        btb_57 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_58 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h3a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_58 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_58 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_58 <= btb_510;
      end else begin
        btb_58 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_59 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h3b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_59 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_59 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_59 <= btb_510;
      end else begin
        btb_59 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_60 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h3c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_60 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_60 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_60 <= btb_510;
      end else begin
        btb_60 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_61 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h3d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_61 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_61 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_61 <= btb_510;
      end else begin
        btb_61 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_62 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h3e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_62 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_62 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_62 <= btb_510;
      end else begin
        btb_62 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_63 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_63 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_63 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_63 <= btb_510;
      end else begin
        btb_63 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_64 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h40 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_64 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_64 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_64 <= btb_510;
      end else begin
        btb_64 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_65 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h41 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_65 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_65 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_65 <= btb_510;
      end else begin
        btb_65 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_66 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h42 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_66 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_66 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_66 <= btb_510;
      end else begin
        btb_66 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_67 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h43 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_67 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_67 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_67 <= btb_510;
      end else begin
        btb_67 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_68 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h44 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_68 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_68 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_68 <= btb_510;
      end else begin
        btb_68 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_69 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h45 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_69 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_69 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_69 <= btb_510;
      end else begin
        btb_69 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_70 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h46 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_70 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_70 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_70 <= btb_510;
      end else begin
        btb_70 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_71 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h47 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_71 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_71 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_71 <= btb_510;
      end else begin
        btb_71 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_72 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h48 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_72 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_72 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_72 <= btb_510;
      end else begin
        btb_72 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_73 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h49 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_73 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_73 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_73 <= btb_510;
      end else begin
        btb_73 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_74 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h4a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_74 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_74 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_74 <= btb_510;
      end else begin
        btb_74 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_75 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h4b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_75 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_75 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_75 <= btb_510;
      end else begin
        btb_75 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_76 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h4c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_76 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_76 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_76 <= btb_510;
      end else begin
        btb_76 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_77 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h4d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_77 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_77 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_77 <= btb_510;
      end else begin
        btb_77 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_78 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h4e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_78 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_78 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_78 <= btb_510;
      end else begin
        btb_78 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_79 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h4f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_79 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_79 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_79 <= btb_510;
      end else begin
        btb_79 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_80 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h50 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_80 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_80 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_80 <= btb_510;
      end else begin
        btb_80 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_81 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h51 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_81 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_81 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_81 <= btb_510;
      end else begin
        btb_81 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_82 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h52 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_82 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_82 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_82 <= btb_510;
      end else begin
        btb_82 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_83 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h53 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_83 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_83 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_83 <= btb_510;
      end else begin
        btb_83 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_84 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h54 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_84 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_84 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_84 <= btb_510;
      end else begin
        btb_84 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_85 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h55 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_85 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_85 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_85 <= btb_510;
      end else begin
        btb_85 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_86 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h56 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_86 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_86 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_86 <= btb_510;
      end else begin
        btb_86 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_87 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h57 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_87 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_87 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_87 <= btb_510;
      end else begin
        btb_87 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_88 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h58 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_88 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_88 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_88 <= btb_510;
      end else begin
        btb_88 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_89 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h59 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_89 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_89 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_89 <= btb_510;
      end else begin
        btb_89 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_90 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h5a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_90 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_90 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_90 <= btb_510;
      end else begin
        btb_90 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_91 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h5b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_91 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_91 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_91 <= btb_510;
      end else begin
        btb_91 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_92 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h5c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_92 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_92 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_92 <= btb_510;
      end else begin
        btb_92 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_93 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h5d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_93 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_93 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_93 <= btb_510;
      end else begin
        btb_93 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_94 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h5e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_94 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_94 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_94 <= btb_510;
      end else begin
        btb_94 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_95 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h5f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_95 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_95 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_95 <= btb_510;
      end else begin
        btb_95 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_96 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h60 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_96 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_96 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_96 <= btb_510;
      end else begin
        btb_96 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_97 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h61 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_97 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_97 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_97 <= btb_510;
      end else begin
        btb_97 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_98 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h62 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_98 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_98 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_98 <= btb_510;
      end else begin
        btb_98 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_99 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h63 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_99 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_99 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_99 <= btb_510;
      end else begin
        btb_99 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_100 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h64 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_100 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_100 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_100 <= btb_510;
      end else begin
        btb_100 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_101 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h65 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_101 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_101 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_101 <= btb_510;
      end else begin
        btb_101 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_102 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h66 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_102 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_102 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_102 <= btb_510;
      end else begin
        btb_102 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_103 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h67 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_103 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_103 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_103 <= btb_510;
      end else begin
        btb_103 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_104 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h68 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_104 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_104 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_104 <= btb_510;
      end else begin
        btb_104 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_105 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h69 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_105 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_105 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_105 <= btb_510;
      end else begin
        btb_105 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_106 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h6a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_106 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_106 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_106 <= btb_510;
      end else begin
        btb_106 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_107 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h6b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_107 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_107 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_107 <= btb_510;
      end else begin
        btb_107 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_108 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h6c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_108 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_108 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_108 <= btb_510;
      end else begin
        btb_108 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_109 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h6d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_109 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_109 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_109 <= btb_510;
      end else begin
        btb_109 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_110 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h6e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_110 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_110 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_110 <= btb_510;
      end else begin
        btb_110 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_111 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h6f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_111 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_111 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_111 <= btb_510;
      end else begin
        btb_111 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_112 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h70 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_112 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_112 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_112 <= btb_510;
      end else begin
        btb_112 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_113 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h71 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_113 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_113 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_113 <= btb_510;
      end else begin
        btb_113 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_114 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h72 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_114 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_114 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_114 <= btb_510;
      end else begin
        btb_114 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_115 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h73 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_115 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_115 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_115 <= btb_510;
      end else begin
        btb_115 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_116 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h74 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_116 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_116 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_116 <= btb_510;
      end else begin
        btb_116 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_117 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h75 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_117 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_117 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_117 <= btb_510;
      end else begin
        btb_117 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_118 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h76 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_118 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_118 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_118 <= btb_510;
      end else begin
        btb_118 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_119 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h77 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_119 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_119 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_119 <= btb_510;
      end else begin
        btb_119 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_120 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h78 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_120 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_120 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_120 <= btb_510;
      end else begin
        btb_120 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_121 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h79 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_121 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_121 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_121 <= btb_510;
      end else begin
        btb_121 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_122 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h7a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_122 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_122 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_122 <= btb_510;
      end else begin
        btb_122 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_123 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h7b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_123 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_123 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_123 <= btb_510;
      end else begin
        btb_123 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_124 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h7c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_124 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_124 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_124 <= btb_510;
      end else begin
        btb_124 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_125 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h7d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_125 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_125 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_125 <= btb_510;
      end else begin
        btb_125 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_126 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h7e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_126 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_126 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_126 <= btb_510;
      end else begin
        btb_126 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_127 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h7f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_127 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_127 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_127 <= btb_510;
      end else begin
        btb_127 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_128 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h80 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_128 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_128 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_128 <= btb_510;
      end else begin
        btb_128 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_129 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h81 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_129 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_129 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_129 <= btb_510;
      end else begin
        btb_129 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_130 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h82 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_130 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_130 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_130 <= btb_510;
      end else begin
        btb_130 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_131 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h83 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_131 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_131 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_131 <= btb_510;
      end else begin
        btb_131 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_132 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h84 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_132 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_132 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_132 <= btb_510;
      end else begin
        btb_132 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_133 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h85 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_133 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_133 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_133 <= btb_510;
      end else begin
        btb_133 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_134 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h86 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_134 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_134 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_134 <= btb_510;
      end else begin
        btb_134 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_135 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h87 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_135 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_135 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_135 <= btb_510;
      end else begin
        btb_135 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_136 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h88 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_136 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_136 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_136 <= btb_510;
      end else begin
        btb_136 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_137 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h89 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_137 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_137 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_137 <= btb_510;
      end else begin
        btb_137 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_138 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h8a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_138 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_138 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_138 <= btb_510;
      end else begin
        btb_138 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_139 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h8b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_139 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_139 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_139 <= btb_510;
      end else begin
        btb_139 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_140 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h8c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_140 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_140 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_140 <= btb_510;
      end else begin
        btb_140 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_141 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h8d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_141 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_141 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_141 <= btb_510;
      end else begin
        btb_141 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_142 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h8e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_142 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_142 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_142 <= btb_510;
      end else begin
        btb_142 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_143 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h8f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_143 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_143 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_143 <= btb_510;
      end else begin
        btb_143 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_144 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h90 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_144 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_144 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_144 <= btb_510;
      end else begin
        btb_144 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_145 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h91 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_145 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_145 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_145 <= btb_510;
      end else begin
        btb_145 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_146 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h92 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_146 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_146 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_146 <= btb_510;
      end else begin
        btb_146 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_147 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h93 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_147 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_147 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_147 <= btb_510;
      end else begin
        btb_147 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_148 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h94 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_148 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_148 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_148 <= btb_510;
      end else begin
        btb_148 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_149 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h95 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_149 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_149 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_149 <= btb_510;
      end else begin
        btb_149 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_150 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h96 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_150 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_150 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_150 <= btb_510;
      end else begin
        btb_150 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_151 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h97 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_151 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_151 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_151 <= btb_510;
      end else begin
        btb_151 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_152 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h98 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_152 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_152 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_152 <= btb_510;
      end else begin
        btb_152 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_153 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h99 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_153 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_153 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_153 <= btb_510;
      end else begin
        btb_153 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_154 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h9a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_154 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_154 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_154 <= btb_510;
      end else begin
        btb_154 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_155 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h9b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_155 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_155 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_155 <= btb_510;
      end else begin
        btb_155 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_156 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h9c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_156 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_156 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_156 <= btb_510;
      end else begin
        btb_156 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_157 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h9d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_157 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_157 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_157 <= btb_510;
      end else begin
        btb_157 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_158 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h9e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_158 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_158 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_158 <= btb_510;
      end else begin
        btb_158 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_159 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h9f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_159 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_159 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_159 <= btb_510;
      end else begin
        btb_159 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_160 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_160 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_160 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_160 <= btb_510;
      end else begin
        btb_160 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_161 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_161 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_161 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_161 <= btb_510;
      end else begin
        btb_161 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_162 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_162 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_162 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_162 <= btb_510;
      end else begin
        btb_162 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_163 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_163 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_163 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_163 <= btb_510;
      end else begin
        btb_163 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_164 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_164 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_164 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_164 <= btb_510;
      end else begin
        btb_164 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_165 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_165 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_165 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_165 <= btb_510;
      end else begin
        btb_165 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_166 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_166 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_166 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_166 <= btb_510;
      end else begin
        btb_166 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_167 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_167 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_167 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_167 <= btb_510;
      end else begin
        btb_167 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_168 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_168 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_168 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_168 <= btb_510;
      end else begin
        btb_168 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_169 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_169 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_169 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_169 <= btb_510;
      end else begin
        btb_169 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_170 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'haa == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_170 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_170 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_170 <= btb_510;
      end else begin
        btb_170 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_171 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hab == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_171 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_171 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_171 <= btb_510;
      end else begin
        btb_171 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_172 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hac == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_172 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_172 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_172 <= btb_510;
      end else begin
        btb_172 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_173 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'had == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_173 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_173 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_173 <= btb_510;
      end else begin
        btb_173 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_174 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hae == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_174 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_174 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_174 <= btb_510;
      end else begin
        btb_174 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_175 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'haf == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_175 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_175 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_175 <= btb_510;
      end else begin
        btb_175 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_176 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_176 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_176 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_176 <= btb_510;
      end else begin
        btb_176 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_177 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_177 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_177 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_177 <= btb_510;
      end else begin
        btb_177 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_178 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_178 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_178 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_178 <= btb_510;
      end else begin
        btb_178 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_179 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_179 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_179 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_179 <= btb_510;
      end else begin
        btb_179 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_180 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_180 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_180 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_180 <= btb_510;
      end else begin
        btb_180 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_181 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_181 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_181 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_181 <= btb_510;
      end else begin
        btb_181 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_182 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_182 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_182 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_182 <= btb_510;
      end else begin
        btb_182 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_183 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_183 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_183 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_183 <= btb_510;
      end else begin
        btb_183 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_184 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_184 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_184 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_184 <= btb_510;
      end else begin
        btb_184 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_185 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_185 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_185 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_185 <= btb_510;
      end else begin
        btb_185 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_186 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hba == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_186 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_186 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_186 <= btb_510;
      end else begin
        btb_186 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_187 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hbb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_187 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_187 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_187 <= btb_510;
      end else begin
        btb_187 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_188 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hbc == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_188 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_188 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_188 <= btb_510;
      end else begin
        btb_188 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_189 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hbd == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_189 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_189 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_189 <= btb_510;
      end else begin
        btb_189 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_190 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hbe == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_190 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_190 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_190 <= btb_510;
      end else begin
        btb_190 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_191 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hbf == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_191 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_191 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_191 <= btb_510;
      end else begin
        btb_191 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_192 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_192 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_192 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_192 <= btb_510;
      end else begin
        btb_192 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_193 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_193 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_193 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_193 <= btb_510;
      end else begin
        btb_193 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_194 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_194 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_194 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_194 <= btb_510;
      end else begin
        btb_194 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_195 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_195 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_195 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_195 <= btb_510;
      end else begin
        btb_195 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_196 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_196 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_196 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_196 <= btb_510;
      end else begin
        btb_196 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_197 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_197 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_197 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_197 <= btb_510;
      end else begin
        btb_197 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_198 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_198 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_198 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_198 <= btb_510;
      end else begin
        btb_198 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_199 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_199 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_199 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_199 <= btb_510;
      end else begin
        btb_199 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_200 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_200 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_200 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_200 <= btb_510;
      end else begin
        btb_200 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_201 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_201 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_201 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_201 <= btb_510;
      end else begin
        btb_201 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_202 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hca == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_202 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_202 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_202 <= btb_510;
      end else begin
        btb_202 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_203 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hcb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_203 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_203 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_203 <= btb_510;
      end else begin
        btb_203 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_204 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hcc == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_204 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_204 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_204 <= btb_510;
      end else begin
        btb_204 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_205 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hcd == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_205 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_205 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_205 <= btb_510;
      end else begin
        btb_205 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_206 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hce == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_206 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_206 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_206 <= btb_510;
      end else begin
        btb_206 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_207 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hcf == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_207 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_207 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_207 <= btb_510;
      end else begin
        btb_207 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_208 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_208 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_208 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_208 <= btb_510;
      end else begin
        btb_208 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_209 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_209 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_209 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_209 <= btb_510;
      end else begin
        btb_209 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_210 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_210 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_210 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_210 <= btb_510;
      end else begin
        btb_210 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_211 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_211 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_211 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_211 <= btb_510;
      end else begin
        btb_211 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_212 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_212 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_212 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_212 <= btb_510;
      end else begin
        btb_212 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_213 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_213 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_213 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_213 <= btb_510;
      end else begin
        btb_213 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_214 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_214 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_214 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_214 <= btb_510;
      end else begin
        btb_214 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_215 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_215 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_215 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_215 <= btb_510;
      end else begin
        btb_215 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_216 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_216 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_216 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_216 <= btb_510;
      end else begin
        btb_216 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_217 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_217 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_217 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_217 <= btb_510;
      end else begin
        btb_217 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_218 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hda == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_218 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_218 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_218 <= btb_510;
      end else begin
        btb_218 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_219 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hdb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_219 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_219 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_219 <= btb_510;
      end else begin
        btb_219 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_220 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hdc == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_220 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_220 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_220 <= btb_510;
      end else begin
        btb_220 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_221 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hdd == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_221 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_221 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_221 <= btb_510;
      end else begin
        btb_221 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_222 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hde == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_222 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_222 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_222 <= btb_510;
      end else begin
        btb_222 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_223 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hdf == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_223 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_223 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_223 <= btb_510;
      end else begin
        btb_223 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_224 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_224 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_224 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_224 <= btb_510;
      end else begin
        btb_224 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_225 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_225 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_225 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_225 <= btb_510;
      end else begin
        btb_225 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_226 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_226 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_226 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_226 <= btb_510;
      end else begin
        btb_226 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_227 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_227 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_227 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_227 <= btb_510;
      end else begin
        btb_227 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_228 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_228 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_228 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_228 <= btb_510;
      end else begin
        btb_228 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_229 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_229 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_229 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_229 <= btb_510;
      end else begin
        btb_229 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_230 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_230 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_230 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_230 <= btb_510;
      end else begin
        btb_230 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_231 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_231 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_231 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_231 <= btb_510;
      end else begin
        btb_231 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_232 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_232 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_232 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_232 <= btb_510;
      end else begin
        btb_232 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_233 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_233 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_233 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_233 <= btb_510;
      end else begin
        btb_233 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_234 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hea == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_234 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_234 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_234 <= btb_510;
      end else begin
        btb_234 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_235 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'heb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_235 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_235 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_235 <= btb_510;
      end else begin
        btb_235 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_236 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hec == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_236 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_236 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_236 <= btb_510;
      end else begin
        btb_236 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_237 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hed == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_237 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_237 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_237 <= btb_510;
      end else begin
        btb_237 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_238 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hee == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_238 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_238 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_238 <= btb_510;
      end else begin
        btb_238 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_239 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hef == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_239 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_239 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_239 <= btb_510;
      end else begin
        btb_239 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_240 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_240 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_240 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_240 <= btb_510;
      end else begin
        btb_240 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_241 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_241 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_241 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_241 <= btb_510;
      end else begin
        btb_241 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_242 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_242 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_242 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_242 <= btb_510;
      end else begin
        btb_242 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_243 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_243 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_243 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_243 <= btb_510;
      end else begin
        btb_243 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_244 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_244 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_244 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_244 <= btb_510;
      end else begin
        btb_244 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_245 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_245 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_245 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_245 <= btb_510;
      end else begin
        btb_245 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_246 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_246 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_246 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_246 <= btb_510;
      end else begin
        btb_246 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_247 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_247 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_247 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_247 <= btb_510;
      end else begin
        btb_247 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_248 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_248 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_248 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_248 <= btb_510;
      end else begin
        btb_248 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_249 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_249 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_249 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_249 <= btb_510;
      end else begin
        btb_249 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_250 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hfa == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_250 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_250 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_250 <= btb_510;
      end else begin
        btb_250 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_251 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hfb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_251 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_251 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_251 <= btb_510;
      end else begin
        btb_251 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_252 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hfc == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_252 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_252 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_252 <= btb_510;
      end else begin
        btb_252 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_253 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hfd == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_253 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_253 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_253 <= btb_510;
      end else begin
        btb_253 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_254 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hfe == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_254 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_254 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_254 <= btb_510;
      end else begin
        btb_254 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_255 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hff == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_255 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_255 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_255 <= btb_510;
      end else begin
        btb_255 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_256 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h100 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_256 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_256 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_256 <= btb_510;
      end else begin
        btb_256 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_257 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h101 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_257 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_257 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_257 <= btb_510;
      end else begin
        btb_257 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_258 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h102 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_258 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_258 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_258 <= btb_510;
      end else begin
        btb_258 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_259 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h103 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_259 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_259 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_259 <= btb_510;
      end else begin
        btb_259 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_260 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h104 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_260 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_260 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_260 <= btb_510;
      end else begin
        btb_260 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_261 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h105 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_261 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_261 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_261 <= btb_510;
      end else begin
        btb_261 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_262 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h106 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_262 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_262 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_262 <= btb_510;
      end else begin
        btb_262 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_263 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h107 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_263 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_263 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_263 <= btb_510;
      end else begin
        btb_263 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_264 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h108 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_264 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_264 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_264 <= btb_510;
      end else begin
        btb_264 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_265 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h109 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_265 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_265 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_265 <= btb_510;
      end else begin
        btb_265 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_266 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h10a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_266 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_266 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_266 <= btb_510;
      end else begin
        btb_266 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_267 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h10b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_267 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_267 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_267 <= btb_510;
      end else begin
        btb_267 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_268 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h10c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_268 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_268 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_268 <= btb_510;
      end else begin
        btb_268 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_269 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h10d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_269 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_269 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_269 <= btb_510;
      end else begin
        btb_269 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_270 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h10e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_270 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_270 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_270 <= btb_510;
      end else begin
        btb_270 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_271 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h10f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_271 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_271 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_271 <= btb_510;
      end else begin
        btb_271 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_272 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h110 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_272 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_272 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_272 <= btb_510;
      end else begin
        btb_272 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_273 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h111 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_273 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_273 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_273 <= btb_510;
      end else begin
        btb_273 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_274 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h112 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_274 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_274 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_274 <= btb_510;
      end else begin
        btb_274 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_275 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h113 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_275 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_275 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_275 <= btb_510;
      end else begin
        btb_275 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_276 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h114 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_276 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_276 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_276 <= btb_510;
      end else begin
        btb_276 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_277 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h115 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_277 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_277 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_277 <= btb_510;
      end else begin
        btb_277 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_278 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h116 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_278 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_278 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_278 <= btb_510;
      end else begin
        btb_278 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_279 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h117 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_279 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_279 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_279 <= btb_510;
      end else begin
        btb_279 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_280 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h118 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_280 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_280 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_280 <= btb_510;
      end else begin
        btb_280 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_281 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h119 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_281 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_281 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_281 <= btb_510;
      end else begin
        btb_281 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_282 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h11a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_282 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_282 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_282 <= btb_510;
      end else begin
        btb_282 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_283 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h11b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_283 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_283 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_283 <= btb_510;
      end else begin
        btb_283 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_284 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h11c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_284 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_284 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_284 <= btb_510;
      end else begin
        btb_284 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_285 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h11d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_285 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_285 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_285 <= btb_510;
      end else begin
        btb_285 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_286 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h11e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_286 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_286 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_286 <= btb_510;
      end else begin
        btb_286 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_287 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h11f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_287 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_287 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_287 <= btb_510;
      end else begin
        btb_287 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_288 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h120 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_288 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_288 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_288 <= btb_510;
      end else begin
        btb_288 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_289 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h121 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_289 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_289 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_289 <= btb_510;
      end else begin
        btb_289 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_290 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h122 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_290 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_290 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_290 <= btb_510;
      end else begin
        btb_290 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_291 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h123 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_291 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_291 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_291 <= btb_510;
      end else begin
        btb_291 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_292 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h124 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_292 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_292 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_292 <= btb_510;
      end else begin
        btb_292 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_293 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h125 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_293 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_293 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_293 <= btb_510;
      end else begin
        btb_293 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_294 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h126 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_294 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_294 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_294 <= btb_510;
      end else begin
        btb_294 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_295 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h127 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_295 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_295 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_295 <= btb_510;
      end else begin
        btb_295 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_296 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h128 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_296 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_296 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_296 <= btb_510;
      end else begin
        btb_296 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_297 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h129 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_297 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_297 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_297 <= btb_510;
      end else begin
        btb_297 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_298 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h12a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_298 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_298 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_298 <= btb_510;
      end else begin
        btb_298 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_299 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h12b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_299 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_299 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_299 <= btb_510;
      end else begin
        btb_299 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_300 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h12c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_300 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_300 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_300 <= btb_510;
      end else begin
        btb_300 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_301 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h12d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_301 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_301 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_301 <= btb_510;
      end else begin
        btb_301 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_302 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h12e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_302 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_302 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_302 <= btb_510;
      end else begin
        btb_302 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_303 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h12f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_303 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_303 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_303 <= btb_510;
      end else begin
        btb_303 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_304 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h130 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_304 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_304 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_304 <= btb_510;
      end else begin
        btb_304 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_305 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h131 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_305 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_305 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_305 <= btb_510;
      end else begin
        btb_305 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_306 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h132 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_306 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_306 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_306 <= btb_510;
      end else begin
        btb_306 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_307 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h133 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_307 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_307 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_307 <= btb_510;
      end else begin
        btb_307 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_308 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h134 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_308 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_308 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_308 <= btb_510;
      end else begin
        btb_308 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_309 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h135 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_309 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_309 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_309 <= btb_510;
      end else begin
        btb_309 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_310 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h136 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_310 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_310 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_310 <= btb_510;
      end else begin
        btb_310 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_311 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h137 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_311 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_311 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_311 <= btb_510;
      end else begin
        btb_311 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_312 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h138 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_312 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_312 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_312 <= btb_510;
      end else begin
        btb_312 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_313 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h139 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_313 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_313 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_313 <= btb_510;
      end else begin
        btb_313 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_314 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h13a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_314 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_314 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_314 <= btb_510;
      end else begin
        btb_314 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_315 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h13b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_315 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_315 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_315 <= btb_510;
      end else begin
        btb_315 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_316 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h13c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_316 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_316 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_316 <= btb_510;
      end else begin
        btb_316 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_317 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h13d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_317 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_317 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_317 <= btb_510;
      end else begin
        btb_317 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_318 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h13e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_318 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_318 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_318 <= btb_510;
      end else begin
        btb_318 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_319 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h13f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_319 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_319 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_319 <= btb_510;
      end else begin
        btb_319 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_320 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h140 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_320 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_320 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_320 <= btb_510;
      end else begin
        btb_320 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_321 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h141 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_321 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_321 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_321 <= btb_510;
      end else begin
        btb_321 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_322 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h142 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_322 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_322 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_322 <= btb_510;
      end else begin
        btb_322 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_323 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h143 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_323 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_323 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_323 <= btb_510;
      end else begin
        btb_323 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_324 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h144 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_324 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_324 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_324 <= btb_510;
      end else begin
        btb_324 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_325 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h145 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_325 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_325 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_325 <= btb_510;
      end else begin
        btb_325 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_326 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h146 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_326 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_326 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_326 <= btb_510;
      end else begin
        btb_326 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_327 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h147 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_327 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_327 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_327 <= btb_510;
      end else begin
        btb_327 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_328 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h148 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_328 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_328 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_328 <= btb_510;
      end else begin
        btb_328 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_329 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h149 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_329 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_329 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_329 <= btb_510;
      end else begin
        btb_329 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_330 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h14a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_330 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_330 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_330 <= btb_510;
      end else begin
        btb_330 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_331 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h14b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_331 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_331 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_331 <= btb_510;
      end else begin
        btb_331 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_332 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h14c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_332 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_332 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_332 <= btb_510;
      end else begin
        btb_332 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_333 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h14d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_333 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_333 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_333 <= btb_510;
      end else begin
        btb_333 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_334 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h14e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_334 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_334 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_334 <= btb_510;
      end else begin
        btb_334 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_335 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h14f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_335 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_335 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_335 <= btb_510;
      end else begin
        btb_335 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_336 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h150 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_336 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_336 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_336 <= btb_510;
      end else begin
        btb_336 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_337 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h151 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_337 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_337 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_337 <= btb_510;
      end else begin
        btb_337 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_338 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h152 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_338 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_338 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_338 <= btb_510;
      end else begin
        btb_338 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_339 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h153 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_339 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_339 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_339 <= btb_510;
      end else begin
        btb_339 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_340 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h154 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_340 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_340 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_340 <= btb_510;
      end else begin
        btb_340 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_341 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h155 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_341 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_341 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_341 <= btb_510;
      end else begin
        btb_341 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_342 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h156 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_342 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_342 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_342 <= btb_510;
      end else begin
        btb_342 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_343 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h157 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_343 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_343 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_343 <= btb_510;
      end else begin
        btb_343 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_344 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h158 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_344 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_344 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_344 <= btb_510;
      end else begin
        btb_344 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_345 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h159 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_345 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_345 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_345 <= btb_510;
      end else begin
        btb_345 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_346 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h15a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_346 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_346 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_346 <= btb_510;
      end else begin
        btb_346 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_347 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h15b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_347 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_347 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_347 <= btb_510;
      end else begin
        btb_347 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_348 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h15c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_348 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_348 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_348 <= btb_510;
      end else begin
        btb_348 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_349 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h15d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_349 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_349 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_349 <= btb_510;
      end else begin
        btb_349 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_350 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h15e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_350 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_350 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_350 <= btb_510;
      end else begin
        btb_350 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_351 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h15f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_351 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_351 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_351 <= btb_510;
      end else begin
        btb_351 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_352 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h160 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_352 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_352 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_352 <= btb_510;
      end else begin
        btb_352 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_353 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h161 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_353 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_353 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_353 <= btb_510;
      end else begin
        btb_353 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_354 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h162 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_354 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_354 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_354 <= btb_510;
      end else begin
        btb_354 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_355 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h163 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_355 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_355 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_355 <= btb_510;
      end else begin
        btb_355 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_356 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h164 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_356 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_356 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_356 <= btb_510;
      end else begin
        btb_356 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_357 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h165 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_357 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_357 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_357 <= btb_510;
      end else begin
        btb_357 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_358 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h166 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_358 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_358 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_358 <= btb_510;
      end else begin
        btb_358 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_359 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h167 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_359 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_359 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_359 <= btb_510;
      end else begin
        btb_359 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_360 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h168 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_360 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_360 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_360 <= btb_510;
      end else begin
        btb_360 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_361 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h169 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_361 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_361 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_361 <= btb_510;
      end else begin
        btb_361 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_362 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h16a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_362 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_362 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_362 <= btb_510;
      end else begin
        btb_362 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_363 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h16b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_363 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_363 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_363 <= btb_510;
      end else begin
        btb_363 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_364 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h16c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_364 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_364 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_364 <= btb_510;
      end else begin
        btb_364 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_365 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h16d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_365 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_365 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_365 <= btb_510;
      end else begin
        btb_365 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_366 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h16e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_366 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_366 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_366 <= btb_510;
      end else begin
        btb_366 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_367 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h16f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_367 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_367 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_367 <= btb_510;
      end else begin
        btb_367 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_368 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h170 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_368 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_368 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_368 <= btb_510;
      end else begin
        btb_368 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_369 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h171 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_369 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_369 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_369 <= btb_510;
      end else begin
        btb_369 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_370 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h172 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_370 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_370 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_370 <= btb_510;
      end else begin
        btb_370 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_371 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h173 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_371 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_371 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_371 <= btb_510;
      end else begin
        btb_371 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_372 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h174 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_372 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_372 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_372 <= btb_510;
      end else begin
        btb_372 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_373 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h175 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_373 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_373 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_373 <= btb_510;
      end else begin
        btb_373 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_374 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h176 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_374 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_374 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_374 <= btb_510;
      end else begin
        btb_374 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_375 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h177 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_375 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_375 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_375 <= btb_510;
      end else begin
        btb_375 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_376 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h178 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_376 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_376 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_376 <= btb_510;
      end else begin
        btb_376 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_377 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h179 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_377 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_377 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_377 <= btb_510;
      end else begin
        btb_377 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_378 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h17a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_378 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_378 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_378 <= btb_510;
      end else begin
        btb_378 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_379 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h17b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_379 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_379 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_379 <= btb_510;
      end else begin
        btb_379 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_380 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h17c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_380 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_380 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_380 <= btb_510;
      end else begin
        btb_380 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_381 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h17d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_381 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_381 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_381 <= btb_510;
      end else begin
        btb_381 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_382 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h17e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_382 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_382 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_382 <= btb_510;
      end else begin
        btb_382 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_383 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h17f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_383 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_383 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_383 <= btb_510;
      end else begin
        btb_383 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_384 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h180 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_384 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_384 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_384 <= btb_510;
      end else begin
        btb_384 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_385 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h181 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_385 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_385 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_385 <= btb_510;
      end else begin
        btb_385 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_386 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h182 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_386 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_386 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_386 <= btb_510;
      end else begin
        btb_386 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_387 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h183 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_387 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_387 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_387 <= btb_510;
      end else begin
        btb_387 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_388 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h184 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_388 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_388 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_388 <= btb_510;
      end else begin
        btb_388 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_389 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h185 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_389 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_389 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_389 <= btb_510;
      end else begin
        btb_389 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_390 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h186 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_390 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_390 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_390 <= btb_510;
      end else begin
        btb_390 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_391 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h187 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_391 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_391 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_391 <= btb_510;
      end else begin
        btb_391 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_392 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h188 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_392 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_392 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_392 <= btb_510;
      end else begin
        btb_392 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_393 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h189 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_393 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_393 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_393 <= btb_510;
      end else begin
        btb_393 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_394 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h18a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_394 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_394 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_394 <= btb_510;
      end else begin
        btb_394 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_395 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h18b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_395 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_395 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_395 <= btb_510;
      end else begin
        btb_395 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_396 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h18c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_396 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_396 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_396 <= btb_510;
      end else begin
        btb_396 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_397 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h18d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_397 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_397 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_397 <= btb_510;
      end else begin
        btb_397 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_398 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h18e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_398 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_398 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_398 <= btb_510;
      end else begin
        btb_398 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_399 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h18f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_399 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_399 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_399 <= btb_510;
      end else begin
        btb_399 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_400 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h190 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_400 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_400 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_400 <= btb_510;
      end else begin
        btb_400 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_401 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h191 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_401 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_401 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_401 <= btb_510;
      end else begin
        btb_401 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_402 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h192 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_402 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_402 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_402 <= btb_510;
      end else begin
        btb_402 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_403 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h193 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_403 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_403 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_403 <= btb_510;
      end else begin
        btb_403 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_404 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h194 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_404 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_404 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_404 <= btb_510;
      end else begin
        btb_404 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_405 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h195 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_405 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_405 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_405 <= btb_510;
      end else begin
        btb_405 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_406 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h196 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_406 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_406 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_406 <= btb_510;
      end else begin
        btb_406 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_407 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h197 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_407 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_407 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_407 <= btb_510;
      end else begin
        btb_407 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_408 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h198 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_408 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_408 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_408 <= btb_510;
      end else begin
        btb_408 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_409 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h199 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_409 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_409 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_409 <= btb_510;
      end else begin
        btb_409 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_410 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h19a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_410 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_410 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_410 <= btb_510;
      end else begin
        btb_410 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_411 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h19b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_411 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_411 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_411 <= btb_510;
      end else begin
        btb_411 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_412 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h19c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_412 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_412 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_412 <= btb_510;
      end else begin
        btb_412 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_413 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h19d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_413 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_413 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_413 <= btb_510;
      end else begin
        btb_413 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_414 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h19e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_414 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_414 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_414 <= btb_510;
      end else begin
        btb_414 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_415 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h19f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_415 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_415 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_415 <= btb_510;
      end else begin
        btb_415 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_416 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_416 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_416 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_416 <= btb_510;
      end else begin
        btb_416 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_417 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_417 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_417 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_417 <= btb_510;
      end else begin
        btb_417 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_418 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_418 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_418 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_418 <= btb_510;
      end else begin
        btb_418 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_419 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_419 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_419 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_419 <= btb_510;
      end else begin
        btb_419 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_420 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_420 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_420 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_420 <= btb_510;
      end else begin
        btb_420 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_421 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_421 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_421 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_421 <= btb_510;
      end else begin
        btb_421 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_422 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_422 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_422 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_422 <= btb_510;
      end else begin
        btb_422 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_423 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_423 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_423 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_423 <= btb_510;
      end else begin
        btb_423 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_424 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_424 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_424 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_424 <= btb_510;
      end else begin
        btb_424 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_425 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_425 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_425 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_425 <= btb_510;
      end else begin
        btb_425 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_426 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1aa == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_426 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_426 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_426 <= btb_510;
      end else begin
        btb_426 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_427 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ab == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_427 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_427 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_427 <= btb_510;
      end else begin
        btb_427 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_428 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ac == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_428 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_428 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_428 <= btb_510;
      end else begin
        btb_428 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_429 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ad == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_429 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_429 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_429 <= btb_510;
      end else begin
        btb_429 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_430 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ae == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_430 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_430 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_430 <= btb_510;
      end else begin
        btb_430 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_431 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1af == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_431 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_431 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_431 <= btb_510;
      end else begin
        btb_431 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_432 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_432 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_432 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_432 <= btb_510;
      end else begin
        btb_432 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_433 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_433 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_433 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_433 <= btb_510;
      end else begin
        btb_433 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_434 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_434 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_434 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_434 <= btb_510;
      end else begin
        btb_434 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_435 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_435 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_435 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_435 <= btb_510;
      end else begin
        btb_435 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_436 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_436 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_436 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_436 <= btb_510;
      end else begin
        btb_436 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_437 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_437 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_437 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_437 <= btb_510;
      end else begin
        btb_437 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_438 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_438 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_438 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_438 <= btb_510;
      end else begin
        btb_438 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_439 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_439 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_439 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_439 <= btb_510;
      end else begin
        btb_439 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_440 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_440 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_440 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_440 <= btb_510;
      end else begin
        btb_440 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_441 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_441 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_441 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_441 <= btb_510;
      end else begin
        btb_441 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_442 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ba == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_442 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_442 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_442 <= btb_510;
      end else begin
        btb_442 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_443 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1bb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_443 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_443 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_443 <= btb_510;
      end else begin
        btb_443 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_444 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1bc == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_444 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_444 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_444 <= btb_510;
      end else begin
        btb_444 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_445 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1bd == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_445 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_445 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_445 <= btb_510;
      end else begin
        btb_445 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_446 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1be == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_446 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_446 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_446 <= btb_510;
      end else begin
        btb_446 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_447 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1bf == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_447 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_447 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_447 <= btb_510;
      end else begin
        btb_447 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_448 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_448 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_448 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_448 <= btb_510;
      end else begin
        btb_448 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_449 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_449 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_449 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_449 <= btb_510;
      end else begin
        btb_449 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_450 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_450 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_450 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_450 <= btb_510;
      end else begin
        btb_450 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_451 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_451 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_451 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_451 <= btb_510;
      end else begin
        btb_451 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_452 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_452 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_452 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_452 <= btb_510;
      end else begin
        btb_452 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_453 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_453 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_453 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_453 <= btb_510;
      end else begin
        btb_453 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_454 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_454 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_454 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_454 <= btb_510;
      end else begin
        btb_454 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_455 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_455 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_455 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_455 <= btb_510;
      end else begin
        btb_455 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_456 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_456 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_456 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_456 <= btb_510;
      end else begin
        btb_456 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_457 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_457 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_457 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_457 <= btb_510;
      end else begin
        btb_457 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_458 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ca == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_458 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_458 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_458 <= btb_510;
      end else begin
        btb_458 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_459 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1cb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_459 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_459 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_459 <= btb_510;
      end else begin
        btb_459 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_460 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1cc == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_460 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_460 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_460 <= btb_510;
      end else begin
        btb_460 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_461 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1cd == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_461 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_461 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_461 <= btb_510;
      end else begin
        btb_461 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_462 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ce == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_462 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_462 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_462 <= btb_510;
      end else begin
        btb_462 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_463 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1cf == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_463 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_463 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_463 <= btb_510;
      end else begin
        btb_463 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_464 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_464 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_464 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_464 <= btb_510;
      end else begin
        btb_464 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_465 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_465 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_465 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_465 <= btb_510;
      end else begin
        btb_465 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_466 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_466 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_466 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_466 <= btb_510;
      end else begin
        btb_466 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_467 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_467 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_467 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_467 <= btb_510;
      end else begin
        btb_467 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_468 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_468 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_468 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_468 <= btb_510;
      end else begin
        btb_468 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_469 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_469 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_469 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_469 <= btb_510;
      end else begin
        btb_469 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_470 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_470 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_470 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_470 <= btb_510;
      end else begin
        btb_470 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_471 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_471 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_471 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_471 <= btb_510;
      end else begin
        btb_471 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_472 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_472 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_472 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_472 <= btb_510;
      end else begin
        btb_472 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_473 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_473 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_473 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_473 <= btb_510;
      end else begin
        btb_473 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_474 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1da == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_474 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_474 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_474 <= btb_510;
      end else begin
        btb_474 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_475 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1db == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_475 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_475 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_475 <= btb_510;
      end else begin
        btb_475 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_476 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1dc == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_476 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_476 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_476 <= btb_510;
      end else begin
        btb_476 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_477 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1dd == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_477 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_477 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_477 <= btb_510;
      end else begin
        btb_477 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_478 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1de == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_478 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_478 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_478 <= btb_510;
      end else begin
        btb_478 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_479 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1df == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_479 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_479 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_479 <= btb_510;
      end else begin
        btb_479 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_480 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_480 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_480 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_480 <= btb_510;
      end else begin
        btb_480 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_481 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_481 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_481 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_481 <= btb_510;
      end else begin
        btb_481 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_482 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_482 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_482 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_482 <= btb_510;
      end else begin
        btb_482 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_483 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_483 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_483 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_483 <= btb_510;
      end else begin
        btb_483 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_484 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_484 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_484 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_484 <= btb_510;
      end else begin
        btb_484 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_485 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_485 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_485 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_485 <= btb_510;
      end else begin
        btb_485 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_486 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_486 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_486 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_486 <= btb_510;
      end else begin
        btb_486 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_487 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_487 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_487 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_487 <= btb_510;
      end else begin
        btb_487 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_488 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_488 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_488 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_488 <= btb_510;
      end else begin
        btb_488 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_489 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_489 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_489 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_489 <= btb_510;
      end else begin
        btb_489 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_490 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ea == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_490 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_490 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_490 <= btb_510;
      end else begin
        btb_490 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_491 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1eb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_491 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_491 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_491 <= btb_510;
      end else begin
        btb_491 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_492 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ec == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_492 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_492 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_492 <= btb_510;
      end else begin
        btb_492 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_493 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ed == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_493 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_493 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_493 <= btb_510;
      end else begin
        btb_493 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_494 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ee == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_494 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_494 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_494 <= btb_510;
      end else begin
        btb_494 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_495 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ef == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_495 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_495 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_495 <= btb_510;
      end else begin
        btb_495 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_496 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_496 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_496 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_496 <= btb_510;
      end else begin
        btb_496 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_497 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_497 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_497 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_497 <= btb_510;
      end else begin
        btb_497 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_498 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_498 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_498 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_498 <= btb_510;
      end else begin
        btb_498 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_499 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_499 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_499 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_499 <= btb_510;
      end else begin
        btb_499 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_500 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_500 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_500 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_500 <= btb_510;
      end else begin
        btb_500 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_501 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_501 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_501 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_501 <= btb_510;
      end else begin
        btb_501 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_502 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_502 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_502 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_502 <= btb_510;
      end else begin
        btb_502 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_503 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_503 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_503 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_503 <= btb_510;
      end else begin
        btb_503 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_504 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_504 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_504 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_504 <= btb_510;
      end else begin
        btb_504 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_505 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_505 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_505 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_505 <= btb_510;
      end else begin
        btb_505 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_506 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1fa == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_506 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_506 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_506 <= btb_510;
      end else begin
        btb_506 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_507 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1fb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_507 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_507 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_507 <= btb_510;
      end else begin
        btb_507 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_508 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1fc == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_508 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_508 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_508 <= btb_510;
      end else begin
        btb_508 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_509 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1fd == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_509 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_509 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_509 <= btb_510;
      end else begin
        btb_509 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_510 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1fe == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_510 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_510 <= btb_511;
      end else if (!(9'h1fe == io_aw_addr)) begin
        btb_510 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_511 <= 8'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ff == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_511 <= io_in;
      end else if (!(9'h1ff == io_aw_addr)) begin
        if (9'h1fe == io_aw_addr) begin
          btb_511 <= btb_510;
        end else begin
          btb_511 <= _GEN_1021;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  btb_0 = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  btb_1 = _RAND_1[7:0];
  _RAND_2 = {1{`RANDOM}};
  btb_2 = _RAND_2[7:0];
  _RAND_3 = {1{`RANDOM}};
  btb_3 = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  btb_4 = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  btb_5 = _RAND_5[7:0];
  _RAND_6 = {1{`RANDOM}};
  btb_6 = _RAND_6[7:0];
  _RAND_7 = {1{`RANDOM}};
  btb_7 = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  btb_8 = _RAND_8[7:0];
  _RAND_9 = {1{`RANDOM}};
  btb_9 = _RAND_9[7:0];
  _RAND_10 = {1{`RANDOM}};
  btb_10 = _RAND_10[7:0];
  _RAND_11 = {1{`RANDOM}};
  btb_11 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  btb_12 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  btb_13 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  btb_14 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  btb_15 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  btb_16 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  btb_17 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  btb_18 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  btb_19 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  btb_20 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  btb_21 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  btb_22 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  btb_23 = _RAND_23[7:0];
  _RAND_24 = {1{`RANDOM}};
  btb_24 = _RAND_24[7:0];
  _RAND_25 = {1{`RANDOM}};
  btb_25 = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  btb_26 = _RAND_26[7:0];
  _RAND_27 = {1{`RANDOM}};
  btb_27 = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  btb_28 = _RAND_28[7:0];
  _RAND_29 = {1{`RANDOM}};
  btb_29 = _RAND_29[7:0];
  _RAND_30 = {1{`RANDOM}};
  btb_30 = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  btb_31 = _RAND_31[7:0];
  _RAND_32 = {1{`RANDOM}};
  btb_32 = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  btb_33 = _RAND_33[7:0];
  _RAND_34 = {1{`RANDOM}};
  btb_34 = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  btb_35 = _RAND_35[7:0];
  _RAND_36 = {1{`RANDOM}};
  btb_36 = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  btb_37 = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  btb_38 = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  btb_39 = _RAND_39[7:0];
  _RAND_40 = {1{`RANDOM}};
  btb_40 = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  btb_41 = _RAND_41[7:0];
  _RAND_42 = {1{`RANDOM}};
  btb_42 = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  btb_43 = _RAND_43[7:0];
  _RAND_44 = {1{`RANDOM}};
  btb_44 = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  btb_45 = _RAND_45[7:0];
  _RAND_46 = {1{`RANDOM}};
  btb_46 = _RAND_46[7:0];
  _RAND_47 = {1{`RANDOM}};
  btb_47 = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  btb_48 = _RAND_48[7:0];
  _RAND_49 = {1{`RANDOM}};
  btb_49 = _RAND_49[7:0];
  _RAND_50 = {1{`RANDOM}};
  btb_50 = _RAND_50[7:0];
  _RAND_51 = {1{`RANDOM}};
  btb_51 = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  btb_52 = _RAND_52[7:0];
  _RAND_53 = {1{`RANDOM}};
  btb_53 = _RAND_53[7:0];
  _RAND_54 = {1{`RANDOM}};
  btb_54 = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  btb_55 = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  btb_56 = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  btb_57 = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  btb_58 = _RAND_58[7:0];
  _RAND_59 = {1{`RANDOM}};
  btb_59 = _RAND_59[7:0];
  _RAND_60 = {1{`RANDOM}};
  btb_60 = _RAND_60[7:0];
  _RAND_61 = {1{`RANDOM}};
  btb_61 = _RAND_61[7:0];
  _RAND_62 = {1{`RANDOM}};
  btb_62 = _RAND_62[7:0];
  _RAND_63 = {1{`RANDOM}};
  btb_63 = _RAND_63[7:0];
  _RAND_64 = {1{`RANDOM}};
  btb_64 = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  btb_65 = _RAND_65[7:0];
  _RAND_66 = {1{`RANDOM}};
  btb_66 = _RAND_66[7:0];
  _RAND_67 = {1{`RANDOM}};
  btb_67 = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  btb_68 = _RAND_68[7:0];
  _RAND_69 = {1{`RANDOM}};
  btb_69 = _RAND_69[7:0];
  _RAND_70 = {1{`RANDOM}};
  btb_70 = _RAND_70[7:0];
  _RAND_71 = {1{`RANDOM}};
  btb_71 = _RAND_71[7:0];
  _RAND_72 = {1{`RANDOM}};
  btb_72 = _RAND_72[7:0];
  _RAND_73 = {1{`RANDOM}};
  btb_73 = _RAND_73[7:0];
  _RAND_74 = {1{`RANDOM}};
  btb_74 = _RAND_74[7:0];
  _RAND_75 = {1{`RANDOM}};
  btb_75 = _RAND_75[7:0];
  _RAND_76 = {1{`RANDOM}};
  btb_76 = _RAND_76[7:0];
  _RAND_77 = {1{`RANDOM}};
  btb_77 = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  btb_78 = _RAND_78[7:0];
  _RAND_79 = {1{`RANDOM}};
  btb_79 = _RAND_79[7:0];
  _RAND_80 = {1{`RANDOM}};
  btb_80 = _RAND_80[7:0];
  _RAND_81 = {1{`RANDOM}};
  btb_81 = _RAND_81[7:0];
  _RAND_82 = {1{`RANDOM}};
  btb_82 = _RAND_82[7:0];
  _RAND_83 = {1{`RANDOM}};
  btb_83 = _RAND_83[7:0];
  _RAND_84 = {1{`RANDOM}};
  btb_84 = _RAND_84[7:0];
  _RAND_85 = {1{`RANDOM}};
  btb_85 = _RAND_85[7:0];
  _RAND_86 = {1{`RANDOM}};
  btb_86 = _RAND_86[7:0];
  _RAND_87 = {1{`RANDOM}};
  btb_87 = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  btb_88 = _RAND_88[7:0];
  _RAND_89 = {1{`RANDOM}};
  btb_89 = _RAND_89[7:0];
  _RAND_90 = {1{`RANDOM}};
  btb_90 = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  btb_91 = _RAND_91[7:0];
  _RAND_92 = {1{`RANDOM}};
  btb_92 = _RAND_92[7:0];
  _RAND_93 = {1{`RANDOM}};
  btb_93 = _RAND_93[7:0];
  _RAND_94 = {1{`RANDOM}};
  btb_94 = _RAND_94[7:0];
  _RAND_95 = {1{`RANDOM}};
  btb_95 = _RAND_95[7:0];
  _RAND_96 = {1{`RANDOM}};
  btb_96 = _RAND_96[7:0];
  _RAND_97 = {1{`RANDOM}};
  btb_97 = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  btb_98 = _RAND_98[7:0];
  _RAND_99 = {1{`RANDOM}};
  btb_99 = _RAND_99[7:0];
  _RAND_100 = {1{`RANDOM}};
  btb_100 = _RAND_100[7:0];
  _RAND_101 = {1{`RANDOM}};
  btb_101 = _RAND_101[7:0];
  _RAND_102 = {1{`RANDOM}};
  btb_102 = _RAND_102[7:0];
  _RAND_103 = {1{`RANDOM}};
  btb_103 = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  btb_104 = _RAND_104[7:0];
  _RAND_105 = {1{`RANDOM}};
  btb_105 = _RAND_105[7:0];
  _RAND_106 = {1{`RANDOM}};
  btb_106 = _RAND_106[7:0];
  _RAND_107 = {1{`RANDOM}};
  btb_107 = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  btb_108 = _RAND_108[7:0];
  _RAND_109 = {1{`RANDOM}};
  btb_109 = _RAND_109[7:0];
  _RAND_110 = {1{`RANDOM}};
  btb_110 = _RAND_110[7:0];
  _RAND_111 = {1{`RANDOM}};
  btb_111 = _RAND_111[7:0];
  _RAND_112 = {1{`RANDOM}};
  btb_112 = _RAND_112[7:0];
  _RAND_113 = {1{`RANDOM}};
  btb_113 = _RAND_113[7:0];
  _RAND_114 = {1{`RANDOM}};
  btb_114 = _RAND_114[7:0];
  _RAND_115 = {1{`RANDOM}};
  btb_115 = _RAND_115[7:0];
  _RAND_116 = {1{`RANDOM}};
  btb_116 = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  btb_117 = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  btb_118 = _RAND_118[7:0];
  _RAND_119 = {1{`RANDOM}};
  btb_119 = _RAND_119[7:0];
  _RAND_120 = {1{`RANDOM}};
  btb_120 = _RAND_120[7:0];
  _RAND_121 = {1{`RANDOM}};
  btb_121 = _RAND_121[7:0];
  _RAND_122 = {1{`RANDOM}};
  btb_122 = _RAND_122[7:0];
  _RAND_123 = {1{`RANDOM}};
  btb_123 = _RAND_123[7:0];
  _RAND_124 = {1{`RANDOM}};
  btb_124 = _RAND_124[7:0];
  _RAND_125 = {1{`RANDOM}};
  btb_125 = _RAND_125[7:0];
  _RAND_126 = {1{`RANDOM}};
  btb_126 = _RAND_126[7:0];
  _RAND_127 = {1{`RANDOM}};
  btb_127 = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  btb_128 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  btb_129 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  btb_130 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  btb_131 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  btb_132 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  btb_133 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  btb_134 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  btb_135 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  btb_136 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  btb_137 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  btb_138 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  btb_139 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  btb_140 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  btb_141 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  btb_142 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  btb_143 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  btb_144 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  btb_145 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  btb_146 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  btb_147 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  btb_148 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  btb_149 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  btb_150 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  btb_151 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  btb_152 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  btb_153 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  btb_154 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  btb_155 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  btb_156 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  btb_157 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  btb_158 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  btb_159 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  btb_160 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  btb_161 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  btb_162 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  btb_163 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  btb_164 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  btb_165 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  btb_166 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  btb_167 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  btb_168 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  btb_169 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  btb_170 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  btb_171 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  btb_172 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  btb_173 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  btb_174 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  btb_175 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  btb_176 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  btb_177 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  btb_178 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  btb_179 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  btb_180 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  btb_181 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  btb_182 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  btb_183 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  btb_184 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  btb_185 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  btb_186 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  btb_187 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  btb_188 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  btb_189 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  btb_190 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  btb_191 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  btb_192 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  btb_193 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  btb_194 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  btb_195 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  btb_196 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  btb_197 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  btb_198 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  btb_199 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  btb_200 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  btb_201 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  btb_202 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  btb_203 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  btb_204 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  btb_205 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  btb_206 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  btb_207 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  btb_208 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  btb_209 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  btb_210 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  btb_211 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  btb_212 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  btb_213 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  btb_214 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  btb_215 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  btb_216 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  btb_217 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  btb_218 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  btb_219 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  btb_220 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  btb_221 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  btb_222 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  btb_223 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  btb_224 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  btb_225 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  btb_226 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  btb_227 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  btb_228 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  btb_229 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  btb_230 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  btb_231 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  btb_232 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  btb_233 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  btb_234 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  btb_235 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  btb_236 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  btb_237 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  btb_238 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  btb_239 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  btb_240 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  btb_241 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  btb_242 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  btb_243 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  btb_244 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  btb_245 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  btb_246 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  btb_247 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  btb_248 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  btb_249 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  btb_250 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  btb_251 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  btb_252 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  btb_253 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  btb_254 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  btb_255 = _RAND_255[7:0];
  _RAND_256 = {1{`RANDOM}};
  btb_256 = _RAND_256[7:0];
  _RAND_257 = {1{`RANDOM}};
  btb_257 = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  btb_258 = _RAND_258[7:0];
  _RAND_259 = {1{`RANDOM}};
  btb_259 = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  btb_260 = _RAND_260[7:0];
  _RAND_261 = {1{`RANDOM}};
  btb_261 = _RAND_261[7:0];
  _RAND_262 = {1{`RANDOM}};
  btb_262 = _RAND_262[7:0];
  _RAND_263 = {1{`RANDOM}};
  btb_263 = _RAND_263[7:0];
  _RAND_264 = {1{`RANDOM}};
  btb_264 = _RAND_264[7:0];
  _RAND_265 = {1{`RANDOM}};
  btb_265 = _RAND_265[7:0];
  _RAND_266 = {1{`RANDOM}};
  btb_266 = _RAND_266[7:0];
  _RAND_267 = {1{`RANDOM}};
  btb_267 = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  btb_268 = _RAND_268[7:0];
  _RAND_269 = {1{`RANDOM}};
  btb_269 = _RAND_269[7:0];
  _RAND_270 = {1{`RANDOM}};
  btb_270 = _RAND_270[7:0];
  _RAND_271 = {1{`RANDOM}};
  btb_271 = _RAND_271[7:0];
  _RAND_272 = {1{`RANDOM}};
  btb_272 = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  btb_273 = _RAND_273[7:0];
  _RAND_274 = {1{`RANDOM}};
  btb_274 = _RAND_274[7:0];
  _RAND_275 = {1{`RANDOM}};
  btb_275 = _RAND_275[7:0];
  _RAND_276 = {1{`RANDOM}};
  btb_276 = _RAND_276[7:0];
  _RAND_277 = {1{`RANDOM}};
  btb_277 = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  btb_278 = _RAND_278[7:0];
  _RAND_279 = {1{`RANDOM}};
  btb_279 = _RAND_279[7:0];
  _RAND_280 = {1{`RANDOM}};
  btb_280 = _RAND_280[7:0];
  _RAND_281 = {1{`RANDOM}};
  btb_281 = _RAND_281[7:0];
  _RAND_282 = {1{`RANDOM}};
  btb_282 = _RAND_282[7:0];
  _RAND_283 = {1{`RANDOM}};
  btb_283 = _RAND_283[7:0];
  _RAND_284 = {1{`RANDOM}};
  btb_284 = _RAND_284[7:0];
  _RAND_285 = {1{`RANDOM}};
  btb_285 = _RAND_285[7:0];
  _RAND_286 = {1{`RANDOM}};
  btb_286 = _RAND_286[7:0];
  _RAND_287 = {1{`RANDOM}};
  btb_287 = _RAND_287[7:0];
  _RAND_288 = {1{`RANDOM}};
  btb_288 = _RAND_288[7:0];
  _RAND_289 = {1{`RANDOM}};
  btb_289 = _RAND_289[7:0];
  _RAND_290 = {1{`RANDOM}};
  btb_290 = _RAND_290[7:0];
  _RAND_291 = {1{`RANDOM}};
  btb_291 = _RAND_291[7:0];
  _RAND_292 = {1{`RANDOM}};
  btb_292 = _RAND_292[7:0];
  _RAND_293 = {1{`RANDOM}};
  btb_293 = _RAND_293[7:0];
  _RAND_294 = {1{`RANDOM}};
  btb_294 = _RAND_294[7:0];
  _RAND_295 = {1{`RANDOM}};
  btb_295 = _RAND_295[7:0];
  _RAND_296 = {1{`RANDOM}};
  btb_296 = _RAND_296[7:0];
  _RAND_297 = {1{`RANDOM}};
  btb_297 = _RAND_297[7:0];
  _RAND_298 = {1{`RANDOM}};
  btb_298 = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  btb_299 = _RAND_299[7:0];
  _RAND_300 = {1{`RANDOM}};
  btb_300 = _RAND_300[7:0];
  _RAND_301 = {1{`RANDOM}};
  btb_301 = _RAND_301[7:0];
  _RAND_302 = {1{`RANDOM}};
  btb_302 = _RAND_302[7:0];
  _RAND_303 = {1{`RANDOM}};
  btb_303 = _RAND_303[7:0];
  _RAND_304 = {1{`RANDOM}};
  btb_304 = _RAND_304[7:0];
  _RAND_305 = {1{`RANDOM}};
  btb_305 = _RAND_305[7:0];
  _RAND_306 = {1{`RANDOM}};
  btb_306 = _RAND_306[7:0];
  _RAND_307 = {1{`RANDOM}};
  btb_307 = _RAND_307[7:0];
  _RAND_308 = {1{`RANDOM}};
  btb_308 = _RAND_308[7:0];
  _RAND_309 = {1{`RANDOM}};
  btb_309 = _RAND_309[7:0];
  _RAND_310 = {1{`RANDOM}};
  btb_310 = _RAND_310[7:0];
  _RAND_311 = {1{`RANDOM}};
  btb_311 = _RAND_311[7:0];
  _RAND_312 = {1{`RANDOM}};
  btb_312 = _RAND_312[7:0];
  _RAND_313 = {1{`RANDOM}};
  btb_313 = _RAND_313[7:0];
  _RAND_314 = {1{`RANDOM}};
  btb_314 = _RAND_314[7:0];
  _RAND_315 = {1{`RANDOM}};
  btb_315 = _RAND_315[7:0];
  _RAND_316 = {1{`RANDOM}};
  btb_316 = _RAND_316[7:0];
  _RAND_317 = {1{`RANDOM}};
  btb_317 = _RAND_317[7:0];
  _RAND_318 = {1{`RANDOM}};
  btb_318 = _RAND_318[7:0];
  _RAND_319 = {1{`RANDOM}};
  btb_319 = _RAND_319[7:0];
  _RAND_320 = {1{`RANDOM}};
  btb_320 = _RAND_320[7:0];
  _RAND_321 = {1{`RANDOM}};
  btb_321 = _RAND_321[7:0];
  _RAND_322 = {1{`RANDOM}};
  btb_322 = _RAND_322[7:0];
  _RAND_323 = {1{`RANDOM}};
  btb_323 = _RAND_323[7:0];
  _RAND_324 = {1{`RANDOM}};
  btb_324 = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  btb_325 = _RAND_325[7:0];
  _RAND_326 = {1{`RANDOM}};
  btb_326 = _RAND_326[7:0];
  _RAND_327 = {1{`RANDOM}};
  btb_327 = _RAND_327[7:0];
  _RAND_328 = {1{`RANDOM}};
  btb_328 = _RAND_328[7:0];
  _RAND_329 = {1{`RANDOM}};
  btb_329 = _RAND_329[7:0];
  _RAND_330 = {1{`RANDOM}};
  btb_330 = _RAND_330[7:0];
  _RAND_331 = {1{`RANDOM}};
  btb_331 = _RAND_331[7:0];
  _RAND_332 = {1{`RANDOM}};
  btb_332 = _RAND_332[7:0];
  _RAND_333 = {1{`RANDOM}};
  btb_333 = _RAND_333[7:0];
  _RAND_334 = {1{`RANDOM}};
  btb_334 = _RAND_334[7:0];
  _RAND_335 = {1{`RANDOM}};
  btb_335 = _RAND_335[7:0];
  _RAND_336 = {1{`RANDOM}};
  btb_336 = _RAND_336[7:0];
  _RAND_337 = {1{`RANDOM}};
  btb_337 = _RAND_337[7:0];
  _RAND_338 = {1{`RANDOM}};
  btb_338 = _RAND_338[7:0];
  _RAND_339 = {1{`RANDOM}};
  btb_339 = _RAND_339[7:0];
  _RAND_340 = {1{`RANDOM}};
  btb_340 = _RAND_340[7:0];
  _RAND_341 = {1{`RANDOM}};
  btb_341 = _RAND_341[7:0];
  _RAND_342 = {1{`RANDOM}};
  btb_342 = _RAND_342[7:0];
  _RAND_343 = {1{`RANDOM}};
  btb_343 = _RAND_343[7:0];
  _RAND_344 = {1{`RANDOM}};
  btb_344 = _RAND_344[7:0];
  _RAND_345 = {1{`RANDOM}};
  btb_345 = _RAND_345[7:0];
  _RAND_346 = {1{`RANDOM}};
  btb_346 = _RAND_346[7:0];
  _RAND_347 = {1{`RANDOM}};
  btb_347 = _RAND_347[7:0];
  _RAND_348 = {1{`RANDOM}};
  btb_348 = _RAND_348[7:0];
  _RAND_349 = {1{`RANDOM}};
  btb_349 = _RAND_349[7:0];
  _RAND_350 = {1{`RANDOM}};
  btb_350 = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  btb_351 = _RAND_351[7:0];
  _RAND_352 = {1{`RANDOM}};
  btb_352 = _RAND_352[7:0];
  _RAND_353 = {1{`RANDOM}};
  btb_353 = _RAND_353[7:0];
  _RAND_354 = {1{`RANDOM}};
  btb_354 = _RAND_354[7:0];
  _RAND_355 = {1{`RANDOM}};
  btb_355 = _RAND_355[7:0];
  _RAND_356 = {1{`RANDOM}};
  btb_356 = _RAND_356[7:0];
  _RAND_357 = {1{`RANDOM}};
  btb_357 = _RAND_357[7:0];
  _RAND_358 = {1{`RANDOM}};
  btb_358 = _RAND_358[7:0];
  _RAND_359 = {1{`RANDOM}};
  btb_359 = _RAND_359[7:0];
  _RAND_360 = {1{`RANDOM}};
  btb_360 = _RAND_360[7:0];
  _RAND_361 = {1{`RANDOM}};
  btb_361 = _RAND_361[7:0];
  _RAND_362 = {1{`RANDOM}};
  btb_362 = _RAND_362[7:0];
  _RAND_363 = {1{`RANDOM}};
  btb_363 = _RAND_363[7:0];
  _RAND_364 = {1{`RANDOM}};
  btb_364 = _RAND_364[7:0];
  _RAND_365 = {1{`RANDOM}};
  btb_365 = _RAND_365[7:0];
  _RAND_366 = {1{`RANDOM}};
  btb_366 = _RAND_366[7:0];
  _RAND_367 = {1{`RANDOM}};
  btb_367 = _RAND_367[7:0];
  _RAND_368 = {1{`RANDOM}};
  btb_368 = _RAND_368[7:0];
  _RAND_369 = {1{`RANDOM}};
  btb_369 = _RAND_369[7:0];
  _RAND_370 = {1{`RANDOM}};
  btb_370 = _RAND_370[7:0];
  _RAND_371 = {1{`RANDOM}};
  btb_371 = _RAND_371[7:0];
  _RAND_372 = {1{`RANDOM}};
  btb_372 = _RAND_372[7:0];
  _RAND_373 = {1{`RANDOM}};
  btb_373 = _RAND_373[7:0];
  _RAND_374 = {1{`RANDOM}};
  btb_374 = _RAND_374[7:0];
  _RAND_375 = {1{`RANDOM}};
  btb_375 = _RAND_375[7:0];
  _RAND_376 = {1{`RANDOM}};
  btb_376 = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  btb_377 = _RAND_377[7:0];
  _RAND_378 = {1{`RANDOM}};
  btb_378 = _RAND_378[7:0];
  _RAND_379 = {1{`RANDOM}};
  btb_379 = _RAND_379[7:0];
  _RAND_380 = {1{`RANDOM}};
  btb_380 = _RAND_380[7:0];
  _RAND_381 = {1{`RANDOM}};
  btb_381 = _RAND_381[7:0];
  _RAND_382 = {1{`RANDOM}};
  btb_382 = _RAND_382[7:0];
  _RAND_383 = {1{`RANDOM}};
  btb_383 = _RAND_383[7:0];
  _RAND_384 = {1{`RANDOM}};
  btb_384 = _RAND_384[7:0];
  _RAND_385 = {1{`RANDOM}};
  btb_385 = _RAND_385[7:0];
  _RAND_386 = {1{`RANDOM}};
  btb_386 = _RAND_386[7:0];
  _RAND_387 = {1{`RANDOM}};
  btb_387 = _RAND_387[7:0];
  _RAND_388 = {1{`RANDOM}};
  btb_388 = _RAND_388[7:0];
  _RAND_389 = {1{`RANDOM}};
  btb_389 = _RAND_389[7:0];
  _RAND_390 = {1{`RANDOM}};
  btb_390 = _RAND_390[7:0];
  _RAND_391 = {1{`RANDOM}};
  btb_391 = _RAND_391[7:0];
  _RAND_392 = {1{`RANDOM}};
  btb_392 = _RAND_392[7:0];
  _RAND_393 = {1{`RANDOM}};
  btb_393 = _RAND_393[7:0];
  _RAND_394 = {1{`RANDOM}};
  btb_394 = _RAND_394[7:0];
  _RAND_395 = {1{`RANDOM}};
  btb_395 = _RAND_395[7:0];
  _RAND_396 = {1{`RANDOM}};
  btb_396 = _RAND_396[7:0];
  _RAND_397 = {1{`RANDOM}};
  btb_397 = _RAND_397[7:0];
  _RAND_398 = {1{`RANDOM}};
  btb_398 = _RAND_398[7:0];
  _RAND_399 = {1{`RANDOM}};
  btb_399 = _RAND_399[7:0];
  _RAND_400 = {1{`RANDOM}};
  btb_400 = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  btb_401 = _RAND_401[7:0];
  _RAND_402 = {1{`RANDOM}};
  btb_402 = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  btb_403 = _RAND_403[7:0];
  _RAND_404 = {1{`RANDOM}};
  btb_404 = _RAND_404[7:0];
  _RAND_405 = {1{`RANDOM}};
  btb_405 = _RAND_405[7:0];
  _RAND_406 = {1{`RANDOM}};
  btb_406 = _RAND_406[7:0];
  _RAND_407 = {1{`RANDOM}};
  btb_407 = _RAND_407[7:0];
  _RAND_408 = {1{`RANDOM}};
  btb_408 = _RAND_408[7:0];
  _RAND_409 = {1{`RANDOM}};
  btb_409 = _RAND_409[7:0];
  _RAND_410 = {1{`RANDOM}};
  btb_410 = _RAND_410[7:0];
  _RAND_411 = {1{`RANDOM}};
  btb_411 = _RAND_411[7:0];
  _RAND_412 = {1{`RANDOM}};
  btb_412 = _RAND_412[7:0];
  _RAND_413 = {1{`RANDOM}};
  btb_413 = _RAND_413[7:0];
  _RAND_414 = {1{`RANDOM}};
  btb_414 = _RAND_414[7:0];
  _RAND_415 = {1{`RANDOM}};
  btb_415 = _RAND_415[7:0];
  _RAND_416 = {1{`RANDOM}};
  btb_416 = _RAND_416[7:0];
  _RAND_417 = {1{`RANDOM}};
  btb_417 = _RAND_417[7:0];
  _RAND_418 = {1{`RANDOM}};
  btb_418 = _RAND_418[7:0];
  _RAND_419 = {1{`RANDOM}};
  btb_419 = _RAND_419[7:0];
  _RAND_420 = {1{`RANDOM}};
  btb_420 = _RAND_420[7:0];
  _RAND_421 = {1{`RANDOM}};
  btb_421 = _RAND_421[7:0];
  _RAND_422 = {1{`RANDOM}};
  btb_422 = _RAND_422[7:0];
  _RAND_423 = {1{`RANDOM}};
  btb_423 = _RAND_423[7:0];
  _RAND_424 = {1{`RANDOM}};
  btb_424 = _RAND_424[7:0];
  _RAND_425 = {1{`RANDOM}};
  btb_425 = _RAND_425[7:0];
  _RAND_426 = {1{`RANDOM}};
  btb_426 = _RAND_426[7:0];
  _RAND_427 = {1{`RANDOM}};
  btb_427 = _RAND_427[7:0];
  _RAND_428 = {1{`RANDOM}};
  btb_428 = _RAND_428[7:0];
  _RAND_429 = {1{`RANDOM}};
  btb_429 = _RAND_429[7:0];
  _RAND_430 = {1{`RANDOM}};
  btb_430 = _RAND_430[7:0];
  _RAND_431 = {1{`RANDOM}};
  btb_431 = _RAND_431[7:0];
  _RAND_432 = {1{`RANDOM}};
  btb_432 = _RAND_432[7:0];
  _RAND_433 = {1{`RANDOM}};
  btb_433 = _RAND_433[7:0];
  _RAND_434 = {1{`RANDOM}};
  btb_434 = _RAND_434[7:0];
  _RAND_435 = {1{`RANDOM}};
  btb_435 = _RAND_435[7:0];
  _RAND_436 = {1{`RANDOM}};
  btb_436 = _RAND_436[7:0];
  _RAND_437 = {1{`RANDOM}};
  btb_437 = _RAND_437[7:0];
  _RAND_438 = {1{`RANDOM}};
  btb_438 = _RAND_438[7:0];
  _RAND_439 = {1{`RANDOM}};
  btb_439 = _RAND_439[7:0];
  _RAND_440 = {1{`RANDOM}};
  btb_440 = _RAND_440[7:0];
  _RAND_441 = {1{`RANDOM}};
  btb_441 = _RAND_441[7:0];
  _RAND_442 = {1{`RANDOM}};
  btb_442 = _RAND_442[7:0];
  _RAND_443 = {1{`RANDOM}};
  btb_443 = _RAND_443[7:0];
  _RAND_444 = {1{`RANDOM}};
  btb_444 = _RAND_444[7:0];
  _RAND_445 = {1{`RANDOM}};
  btb_445 = _RAND_445[7:0];
  _RAND_446 = {1{`RANDOM}};
  btb_446 = _RAND_446[7:0];
  _RAND_447 = {1{`RANDOM}};
  btb_447 = _RAND_447[7:0];
  _RAND_448 = {1{`RANDOM}};
  btb_448 = _RAND_448[7:0];
  _RAND_449 = {1{`RANDOM}};
  btb_449 = _RAND_449[7:0];
  _RAND_450 = {1{`RANDOM}};
  btb_450 = _RAND_450[7:0];
  _RAND_451 = {1{`RANDOM}};
  btb_451 = _RAND_451[7:0];
  _RAND_452 = {1{`RANDOM}};
  btb_452 = _RAND_452[7:0];
  _RAND_453 = {1{`RANDOM}};
  btb_453 = _RAND_453[7:0];
  _RAND_454 = {1{`RANDOM}};
  btb_454 = _RAND_454[7:0];
  _RAND_455 = {1{`RANDOM}};
  btb_455 = _RAND_455[7:0];
  _RAND_456 = {1{`RANDOM}};
  btb_456 = _RAND_456[7:0];
  _RAND_457 = {1{`RANDOM}};
  btb_457 = _RAND_457[7:0];
  _RAND_458 = {1{`RANDOM}};
  btb_458 = _RAND_458[7:0];
  _RAND_459 = {1{`RANDOM}};
  btb_459 = _RAND_459[7:0];
  _RAND_460 = {1{`RANDOM}};
  btb_460 = _RAND_460[7:0];
  _RAND_461 = {1{`RANDOM}};
  btb_461 = _RAND_461[7:0];
  _RAND_462 = {1{`RANDOM}};
  btb_462 = _RAND_462[7:0];
  _RAND_463 = {1{`RANDOM}};
  btb_463 = _RAND_463[7:0];
  _RAND_464 = {1{`RANDOM}};
  btb_464 = _RAND_464[7:0];
  _RAND_465 = {1{`RANDOM}};
  btb_465 = _RAND_465[7:0];
  _RAND_466 = {1{`RANDOM}};
  btb_466 = _RAND_466[7:0];
  _RAND_467 = {1{`RANDOM}};
  btb_467 = _RAND_467[7:0];
  _RAND_468 = {1{`RANDOM}};
  btb_468 = _RAND_468[7:0];
  _RAND_469 = {1{`RANDOM}};
  btb_469 = _RAND_469[7:0];
  _RAND_470 = {1{`RANDOM}};
  btb_470 = _RAND_470[7:0];
  _RAND_471 = {1{`RANDOM}};
  btb_471 = _RAND_471[7:0];
  _RAND_472 = {1{`RANDOM}};
  btb_472 = _RAND_472[7:0];
  _RAND_473 = {1{`RANDOM}};
  btb_473 = _RAND_473[7:0];
  _RAND_474 = {1{`RANDOM}};
  btb_474 = _RAND_474[7:0];
  _RAND_475 = {1{`RANDOM}};
  btb_475 = _RAND_475[7:0];
  _RAND_476 = {1{`RANDOM}};
  btb_476 = _RAND_476[7:0];
  _RAND_477 = {1{`RANDOM}};
  btb_477 = _RAND_477[7:0];
  _RAND_478 = {1{`RANDOM}};
  btb_478 = _RAND_478[7:0];
  _RAND_479 = {1{`RANDOM}};
  btb_479 = _RAND_479[7:0];
  _RAND_480 = {1{`RANDOM}};
  btb_480 = _RAND_480[7:0];
  _RAND_481 = {1{`RANDOM}};
  btb_481 = _RAND_481[7:0];
  _RAND_482 = {1{`RANDOM}};
  btb_482 = _RAND_482[7:0];
  _RAND_483 = {1{`RANDOM}};
  btb_483 = _RAND_483[7:0];
  _RAND_484 = {1{`RANDOM}};
  btb_484 = _RAND_484[7:0];
  _RAND_485 = {1{`RANDOM}};
  btb_485 = _RAND_485[7:0];
  _RAND_486 = {1{`RANDOM}};
  btb_486 = _RAND_486[7:0];
  _RAND_487 = {1{`RANDOM}};
  btb_487 = _RAND_487[7:0];
  _RAND_488 = {1{`RANDOM}};
  btb_488 = _RAND_488[7:0];
  _RAND_489 = {1{`RANDOM}};
  btb_489 = _RAND_489[7:0];
  _RAND_490 = {1{`RANDOM}};
  btb_490 = _RAND_490[7:0];
  _RAND_491 = {1{`RANDOM}};
  btb_491 = _RAND_491[7:0];
  _RAND_492 = {1{`RANDOM}};
  btb_492 = _RAND_492[7:0];
  _RAND_493 = {1{`RANDOM}};
  btb_493 = _RAND_493[7:0];
  _RAND_494 = {1{`RANDOM}};
  btb_494 = _RAND_494[7:0];
  _RAND_495 = {1{`RANDOM}};
  btb_495 = _RAND_495[7:0];
  _RAND_496 = {1{`RANDOM}};
  btb_496 = _RAND_496[7:0];
  _RAND_497 = {1{`RANDOM}};
  btb_497 = _RAND_497[7:0];
  _RAND_498 = {1{`RANDOM}};
  btb_498 = _RAND_498[7:0];
  _RAND_499 = {1{`RANDOM}};
  btb_499 = _RAND_499[7:0];
  _RAND_500 = {1{`RANDOM}};
  btb_500 = _RAND_500[7:0];
  _RAND_501 = {1{`RANDOM}};
  btb_501 = _RAND_501[7:0];
  _RAND_502 = {1{`RANDOM}};
  btb_502 = _RAND_502[7:0];
  _RAND_503 = {1{`RANDOM}};
  btb_503 = _RAND_503[7:0];
  _RAND_504 = {1{`RANDOM}};
  btb_504 = _RAND_504[7:0];
  _RAND_505 = {1{`RANDOM}};
  btb_505 = _RAND_505[7:0];
  _RAND_506 = {1{`RANDOM}};
  btb_506 = _RAND_506[7:0];
  _RAND_507 = {1{`RANDOM}};
  btb_507 = _RAND_507[7:0];
  _RAND_508 = {1{`RANDOM}};
  btb_508 = _RAND_508[7:0];
  _RAND_509 = {1{`RANDOM}};
  btb_509 = _RAND_509[7:0];
  _RAND_510 = {1{`RANDOM}};
  btb_510 = _RAND_510[7:0];
  _RAND_511 = {1{`RANDOM}};
  btb_511 = _RAND_511[7:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    btb_0 = 8'h0;
  end
  if (reset) begin
    btb_1 = 8'h0;
  end
  if (reset) begin
    btb_2 = 8'h0;
  end
  if (reset) begin
    btb_3 = 8'h0;
  end
  if (reset) begin
    btb_4 = 8'h0;
  end
  if (reset) begin
    btb_5 = 8'h0;
  end
  if (reset) begin
    btb_6 = 8'h0;
  end
  if (reset) begin
    btb_7 = 8'h0;
  end
  if (reset) begin
    btb_8 = 8'h0;
  end
  if (reset) begin
    btb_9 = 8'h0;
  end
  if (reset) begin
    btb_10 = 8'h0;
  end
  if (reset) begin
    btb_11 = 8'h0;
  end
  if (reset) begin
    btb_12 = 8'h0;
  end
  if (reset) begin
    btb_13 = 8'h0;
  end
  if (reset) begin
    btb_14 = 8'h0;
  end
  if (reset) begin
    btb_15 = 8'h0;
  end
  if (reset) begin
    btb_16 = 8'h0;
  end
  if (reset) begin
    btb_17 = 8'h0;
  end
  if (reset) begin
    btb_18 = 8'h0;
  end
  if (reset) begin
    btb_19 = 8'h0;
  end
  if (reset) begin
    btb_20 = 8'h0;
  end
  if (reset) begin
    btb_21 = 8'h0;
  end
  if (reset) begin
    btb_22 = 8'h0;
  end
  if (reset) begin
    btb_23 = 8'h0;
  end
  if (reset) begin
    btb_24 = 8'h0;
  end
  if (reset) begin
    btb_25 = 8'h0;
  end
  if (reset) begin
    btb_26 = 8'h0;
  end
  if (reset) begin
    btb_27 = 8'h0;
  end
  if (reset) begin
    btb_28 = 8'h0;
  end
  if (reset) begin
    btb_29 = 8'h0;
  end
  if (reset) begin
    btb_30 = 8'h0;
  end
  if (reset) begin
    btb_31 = 8'h0;
  end
  if (reset) begin
    btb_32 = 8'h0;
  end
  if (reset) begin
    btb_33 = 8'h0;
  end
  if (reset) begin
    btb_34 = 8'h0;
  end
  if (reset) begin
    btb_35 = 8'h0;
  end
  if (reset) begin
    btb_36 = 8'h0;
  end
  if (reset) begin
    btb_37 = 8'h0;
  end
  if (reset) begin
    btb_38 = 8'h0;
  end
  if (reset) begin
    btb_39 = 8'h0;
  end
  if (reset) begin
    btb_40 = 8'h0;
  end
  if (reset) begin
    btb_41 = 8'h0;
  end
  if (reset) begin
    btb_42 = 8'h0;
  end
  if (reset) begin
    btb_43 = 8'h0;
  end
  if (reset) begin
    btb_44 = 8'h0;
  end
  if (reset) begin
    btb_45 = 8'h0;
  end
  if (reset) begin
    btb_46 = 8'h0;
  end
  if (reset) begin
    btb_47 = 8'h0;
  end
  if (reset) begin
    btb_48 = 8'h0;
  end
  if (reset) begin
    btb_49 = 8'h0;
  end
  if (reset) begin
    btb_50 = 8'h0;
  end
  if (reset) begin
    btb_51 = 8'h0;
  end
  if (reset) begin
    btb_52 = 8'h0;
  end
  if (reset) begin
    btb_53 = 8'h0;
  end
  if (reset) begin
    btb_54 = 8'h0;
  end
  if (reset) begin
    btb_55 = 8'h0;
  end
  if (reset) begin
    btb_56 = 8'h0;
  end
  if (reset) begin
    btb_57 = 8'h0;
  end
  if (reset) begin
    btb_58 = 8'h0;
  end
  if (reset) begin
    btb_59 = 8'h0;
  end
  if (reset) begin
    btb_60 = 8'h0;
  end
  if (reset) begin
    btb_61 = 8'h0;
  end
  if (reset) begin
    btb_62 = 8'h0;
  end
  if (reset) begin
    btb_63 = 8'h0;
  end
  if (reset) begin
    btb_64 = 8'h0;
  end
  if (reset) begin
    btb_65 = 8'h0;
  end
  if (reset) begin
    btb_66 = 8'h0;
  end
  if (reset) begin
    btb_67 = 8'h0;
  end
  if (reset) begin
    btb_68 = 8'h0;
  end
  if (reset) begin
    btb_69 = 8'h0;
  end
  if (reset) begin
    btb_70 = 8'h0;
  end
  if (reset) begin
    btb_71 = 8'h0;
  end
  if (reset) begin
    btb_72 = 8'h0;
  end
  if (reset) begin
    btb_73 = 8'h0;
  end
  if (reset) begin
    btb_74 = 8'h0;
  end
  if (reset) begin
    btb_75 = 8'h0;
  end
  if (reset) begin
    btb_76 = 8'h0;
  end
  if (reset) begin
    btb_77 = 8'h0;
  end
  if (reset) begin
    btb_78 = 8'h0;
  end
  if (reset) begin
    btb_79 = 8'h0;
  end
  if (reset) begin
    btb_80 = 8'h0;
  end
  if (reset) begin
    btb_81 = 8'h0;
  end
  if (reset) begin
    btb_82 = 8'h0;
  end
  if (reset) begin
    btb_83 = 8'h0;
  end
  if (reset) begin
    btb_84 = 8'h0;
  end
  if (reset) begin
    btb_85 = 8'h0;
  end
  if (reset) begin
    btb_86 = 8'h0;
  end
  if (reset) begin
    btb_87 = 8'h0;
  end
  if (reset) begin
    btb_88 = 8'h0;
  end
  if (reset) begin
    btb_89 = 8'h0;
  end
  if (reset) begin
    btb_90 = 8'h0;
  end
  if (reset) begin
    btb_91 = 8'h0;
  end
  if (reset) begin
    btb_92 = 8'h0;
  end
  if (reset) begin
    btb_93 = 8'h0;
  end
  if (reset) begin
    btb_94 = 8'h0;
  end
  if (reset) begin
    btb_95 = 8'h0;
  end
  if (reset) begin
    btb_96 = 8'h0;
  end
  if (reset) begin
    btb_97 = 8'h0;
  end
  if (reset) begin
    btb_98 = 8'h0;
  end
  if (reset) begin
    btb_99 = 8'h0;
  end
  if (reset) begin
    btb_100 = 8'h0;
  end
  if (reset) begin
    btb_101 = 8'h0;
  end
  if (reset) begin
    btb_102 = 8'h0;
  end
  if (reset) begin
    btb_103 = 8'h0;
  end
  if (reset) begin
    btb_104 = 8'h0;
  end
  if (reset) begin
    btb_105 = 8'h0;
  end
  if (reset) begin
    btb_106 = 8'h0;
  end
  if (reset) begin
    btb_107 = 8'h0;
  end
  if (reset) begin
    btb_108 = 8'h0;
  end
  if (reset) begin
    btb_109 = 8'h0;
  end
  if (reset) begin
    btb_110 = 8'h0;
  end
  if (reset) begin
    btb_111 = 8'h0;
  end
  if (reset) begin
    btb_112 = 8'h0;
  end
  if (reset) begin
    btb_113 = 8'h0;
  end
  if (reset) begin
    btb_114 = 8'h0;
  end
  if (reset) begin
    btb_115 = 8'h0;
  end
  if (reset) begin
    btb_116 = 8'h0;
  end
  if (reset) begin
    btb_117 = 8'h0;
  end
  if (reset) begin
    btb_118 = 8'h0;
  end
  if (reset) begin
    btb_119 = 8'h0;
  end
  if (reset) begin
    btb_120 = 8'h0;
  end
  if (reset) begin
    btb_121 = 8'h0;
  end
  if (reset) begin
    btb_122 = 8'h0;
  end
  if (reset) begin
    btb_123 = 8'h0;
  end
  if (reset) begin
    btb_124 = 8'h0;
  end
  if (reset) begin
    btb_125 = 8'h0;
  end
  if (reset) begin
    btb_126 = 8'h0;
  end
  if (reset) begin
    btb_127 = 8'h0;
  end
  if (reset) begin
    btb_128 = 8'h0;
  end
  if (reset) begin
    btb_129 = 8'h0;
  end
  if (reset) begin
    btb_130 = 8'h0;
  end
  if (reset) begin
    btb_131 = 8'h0;
  end
  if (reset) begin
    btb_132 = 8'h0;
  end
  if (reset) begin
    btb_133 = 8'h0;
  end
  if (reset) begin
    btb_134 = 8'h0;
  end
  if (reset) begin
    btb_135 = 8'h0;
  end
  if (reset) begin
    btb_136 = 8'h0;
  end
  if (reset) begin
    btb_137 = 8'h0;
  end
  if (reset) begin
    btb_138 = 8'h0;
  end
  if (reset) begin
    btb_139 = 8'h0;
  end
  if (reset) begin
    btb_140 = 8'h0;
  end
  if (reset) begin
    btb_141 = 8'h0;
  end
  if (reset) begin
    btb_142 = 8'h0;
  end
  if (reset) begin
    btb_143 = 8'h0;
  end
  if (reset) begin
    btb_144 = 8'h0;
  end
  if (reset) begin
    btb_145 = 8'h0;
  end
  if (reset) begin
    btb_146 = 8'h0;
  end
  if (reset) begin
    btb_147 = 8'h0;
  end
  if (reset) begin
    btb_148 = 8'h0;
  end
  if (reset) begin
    btb_149 = 8'h0;
  end
  if (reset) begin
    btb_150 = 8'h0;
  end
  if (reset) begin
    btb_151 = 8'h0;
  end
  if (reset) begin
    btb_152 = 8'h0;
  end
  if (reset) begin
    btb_153 = 8'h0;
  end
  if (reset) begin
    btb_154 = 8'h0;
  end
  if (reset) begin
    btb_155 = 8'h0;
  end
  if (reset) begin
    btb_156 = 8'h0;
  end
  if (reset) begin
    btb_157 = 8'h0;
  end
  if (reset) begin
    btb_158 = 8'h0;
  end
  if (reset) begin
    btb_159 = 8'h0;
  end
  if (reset) begin
    btb_160 = 8'h0;
  end
  if (reset) begin
    btb_161 = 8'h0;
  end
  if (reset) begin
    btb_162 = 8'h0;
  end
  if (reset) begin
    btb_163 = 8'h0;
  end
  if (reset) begin
    btb_164 = 8'h0;
  end
  if (reset) begin
    btb_165 = 8'h0;
  end
  if (reset) begin
    btb_166 = 8'h0;
  end
  if (reset) begin
    btb_167 = 8'h0;
  end
  if (reset) begin
    btb_168 = 8'h0;
  end
  if (reset) begin
    btb_169 = 8'h0;
  end
  if (reset) begin
    btb_170 = 8'h0;
  end
  if (reset) begin
    btb_171 = 8'h0;
  end
  if (reset) begin
    btb_172 = 8'h0;
  end
  if (reset) begin
    btb_173 = 8'h0;
  end
  if (reset) begin
    btb_174 = 8'h0;
  end
  if (reset) begin
    btb_175 = 8'h0;
  end
  if (reset) begin
    btb_176 = 8'h0;
  end
  if (reset) begin
    btb_177 = 8'h0;
  end
  if (reset) begin
    btb_178 = 8'h0;
  end
  if (reset) begin
    btb_179 = 8'h0;
  end
  if (reset) begin
    btb_180 = 8'h0;
  end
  if (reset) begin
    btb_181 = 8'h0;
  end
  if (reset) begin
    btb_182 = 8'h0;
  end
  if (reset) begin
    btb_183 = 8'h0;
  end
  if (reset) begin
    btb_184 = 8'h0;
  end
  if (reset) begin
    btb_185 = 8'h0;
  end
  if (reset) begin
    btb_186 = 8'h0;
  end
  if (reset) begin
    btb_187 = 8'h0;
  end
  if (reset) begin
    btb_188 = 8'h0;
  end
  if (reset) begin
    btb_189 = 8'h0;
  end
  if (reset) begin
    btb_190 = 8'h0;
  end
  if (reset) begin
    btb_191 = 8'h0;
  end
  if (reset) begin
    btb_192 = 8'h0;
  end
  if (reset) begin
    btb_193 = 8'h0;
  end
  if (reset) begin
    btb_194 = 8'h0;
  end
  if (reset) begin
    btb_195 = 8'h0;
  end
  if (reset) begin
    btb_196 = 8'h0;
  end
  if (reset) begin
    btb_197 = 8'h0;
  end
  if (reset) begin
    btb_198 = 8'h0;
  end
  if (reset) begin
    btb_199 = 8'h0;
  end
  if (reset) begin
    btb_200 = 8'h0;
  end
  if (reset) begin
    btb_201 = 8'h0;
  end
  if (reset) begin
    btb_202 = 8'h0;
  end
  if (reset) begin
    btb_203 = 8'h0;
  end
  if (reset) begin
    btb_204 = 8'h0;
  end
  if (reset) begin
    btb_205 = 8'h0;
  end
  if (reset) begin
    btb_206 = 8'h0;
  end
  if (reset) begin
    btb_207 = 8'h0;
  end
  if (reset) begin
    btb_208 = 8'h0;
  end
  if (reset) begin
    btb_209 = 8'h0;
  end
  if (reset) begin
    btb_210 = 8'h0;
  end
  if (reset) begin
    btb_211 = 8'h0;
  end
  if (reset) begin
    btb_212 = 8'h0;
  end
  if (reset) begin
    btb_213 = 8'h0;
  end
  if (reset) begin
    btb_214 = 8'h0;
  end
  if (reset) begin
    btb_215 = 8'h0;
  end
  if (reset) begin
    btb_216 = 8'h0;
  end
  if (reset) begin
    btb_217 = 8'h0;
  end
  if (reset) begin
    btb_218 = 8'h0;
  end
  if (reset) begin
    btb_219 = 8'h0;
  end
  if (reset) begin
    btb_220 = 8'h0;
  end
  if (reset) begin
    btb_221 = 8'h0;
  end
  if (reset) begin
    btb_222 = 8'h0;
  end
  if (reset) begin
    btb_223 = 8'h0;
  end
  if (reset) begin
    btb_224 = 8'h0;
  end
  if (reset) begin
    btb_225 = 8'h0;
  end
  if (reset) begin
    btb_226 = 8'h0;
  end
  if (reset) begin
    btb_227 = 8'h0;
  end
  if (reset) begin
    btb_228 = 8'h0;
  end
  if (reset) begin
    btb_229 = 8'h0;
  end
  if (reset) begin
    btb_230 = 8'h0;
  end
  if (reset) begin
    btb_231 = 8'h0;
  end
  if (reset) begin
    btb_232 = 8'h0;
  end
  if (reset) begin
    btb_233 = 8'h0;
  end
  if (reset) begin
    btb_234 = 8'h0;
  end
  if (reset) begin
    btb_235 = 8'h0;
  end
  if (reset) begin
    btb_236 = 8'h0;
  end
  if (reset) begin
    btb_237 = 8'h0;
  end
  if (reset) begin
    btb_238 = 8'h0;
  end
  if (reset) begin
    btb_239 = 8'h0;
  end
  if (reset) begin
    btb_240 = 8'h0;
  end
  if (reset) begin
    btb_241 = 8'h0;
  end
  if (reset) begin
    btb_242 = 8'h0;
  end
  if (reset) begin
    btb_243 = 8'h0;
  end
  if (reset) begin
    btb_244 = 8'h0;
  end
  if (reset) begin
    btb_245 = 8'h0;
  end
  if (reset) begin
    btb_246 = 8'h0;
  end
  if (reset) begin
    btb_247 = 8'h0;
  end
  if (reset) begin
    btb_248 = 8'h0;
  end
  if (reset) begin
    btb_249 = 8'h0;
  end
  if (reset) begin
    btb_250 = 8'h0;
  end
  if (reset) begin
    btb_251 = 8'h0;
  end
  if (reset) begin
    btb_252 = 8'h0;
  end
  if (reset) begin
    btb_253 = 8'h0;
  end
  if (reset) begin
    btb_254 = 8'h0;
  end
  if (reset) begin
    btb_255 = 8'h0;
  end
  if (reset) begin
    btb_256 = 8'h0;
  end
  if (reset) begin
    btb_257 = 8'h0;
  end
  if (reset) begin
    btb_258 = 8'h0;
  end
  if (reset) begin
    btb_259 = 8'h0;
  end
  if (reset) begin
    btb_260 = 8'h0;
  end
  if (reset) begin
    btb_261 = 8'h0;
  end
  if (reset) begin
    btb_262 = 8'h0;
  end
  if (reset) begin
    btb_263 = 8'h0;
  end
  if (reset) begin
    btb_264 = 8'h0;
  end
  if (reset) begin
    btb_265 = 8'h0;
  end
  if (reset) begin
    btb_266 = 8'h0;
  end
  if (reset) begin
    btb_267 = 8'h0;
  end
  if (reset) begin
    btb_268 = 8'h0;
  end
  if (reset) begin
    btb_269 = 8'h0;
  end
  if (reset) begin
    btb_270 = 8'h0;
  end
  if (reset) begin
    btb_271 = 8'h0;
  end
  if (reset) begin
    btb_272 = 8'h0;
  end
  if (reset) begin
    btb_273 = 8'h0;
  end
  if (reset) begin
    btb_274 = 8'h0;
  end
  if (reset) begin
    btb_275 = 8'h0;
  end
  if (reset) begin
    btb_276 = 8'h0;
  end
  if (reset) begin
    btb_277 = 8'h0;
  end
  if (reset) begin
    btb_278 = 8'h0;
  end
  if (reset) begin
    btb_279 = 8'h0;
  end
  if (reset) begin
    btb_280 = 8'h0;
  end
  if (reset) begin
    btb_281 = 8'h0;
  end
  if (reset) begin
    btb_282 = 8'h0;
  end
  if (reset) begin
    btb_283 = 8'h0;
  end
  if (reset) begin
    btb_284 = 8'h0;
  end
  if (reset) begin
    btb_285 = 8'h0;
  end
  if (reset) begin
    btb_286 = 8'h0;
  end
  if (reset) begin
    btb_287 = 8'h0;
  end
  if (reset) begin
    btb_288 = 8'h0;
  end
  if (reset) begin
    btb_289 = 8'h0;
  end
  if (reset) begin
    btb_290 = 8'h0;
  end
  if (reset) begin
    btb_291 = 8'h0;
  end
  if (reset) begin
    btb_292 = 8'h0;
  end
  if (reset) begin
    btb_293 = 8'h0;
  end
  if (reset) begin
    btb_294 = 8'h0;
  end
  if (reset) begin
    btb_295 = 8'h0;
  end
  if (reset) begin
    btb_296 = 8'h0;
  end
  if (reset) begin
    btb_297 = 8'h0;
  end
  if (reset) begin
    btb_298 = 8'h0;
  end
  if (reset) begin
    btb_299 = 8'h0;
  end
  if (reset) begin
    btb_300 = 8'h0;
  end
  if (reset) begin
    btb_301 = 8'h0;
  end
  if (reset) begin
    btb_302 = 8'h0;
  end
  if (reset) begin
    btb_303 = 8'h0;
  end
  if (reset) begin
    btb_304 = 8'h0;
  end
  if (reset) begin
    btb_305 = 8'h0;
  end
  if (reset) begin
    btb_306 = 8'h0;
  end
  if (reset) begin
    btb_307 = 8'h0;
  end
  if (reset) begin
    btb_308 = 8'h0;
  end
  if (reset) begin
    btb_309 = 8'h0;
  end
  if (reset) begin
    btb_310 = 8'h0;
  end
  if (reset) begin
    btb_311 = 8'h0;
  end
  if (reset) begin
    btb_312 = 8'h0;
  end
  if (reset) begin
    btb_313 = 8'h0;
  end
  if (reset) begin
    btb_314 = 8'h0;
  end
  if (reset) begin
    btb_315 = 8'h0;
  end
  if (reset) begin
    btb_316 = 8'h0;
  end
  if (reset) begin
    btb_317 = 8'h0;
  end
  if (reset) begin
    btb_318 = 8'h0;
  end
  if (reset) begin
    btb_319 = 8'h0;
  end
  if (reset) begin
    btb_320 = 8'h0;
  end
  if (reset) begin
    btb_321 = 8'h0;
  end
  if (reset) begin
    btb_322 = 8'h0;
  end
  if (reset) begin
    btb_323 = 8'h0;
  end
  if (reset) begin
    btb_324 = 8'h0;
  end
  if (reset) begin
    btb_325 = 8'h0;
  end
  if (reset) begin
    btb_326 = 8'h0;
  end
  if (reset) begin
    btb_327 = 8'h0;
  end
  if (reset) begin
    btb_328 = 8'h0;
  end
  if (reset) begin
    btb_329 = 8'h0;
  end
  if (reset) begin
    btb_330 = 8'h0;
  end
  if (reset) begin
    btb_331 = 8'h0;
  end
  if (reset) begin
    btb_332 = 8'h0;
  end
  if (reset) begin
    btb_333 = 8'h0;
  end
  if (reset) begin
    btb_334 = 8'h0;
  end
  if (reset) begin
    btb_335 = 8'h0;
  end
  if (reset) begin
    btb_336 = 8'h0;
  end
  if (reset) begin
    btb_337 = 8'h0;
  end
  if (reset) begin
    btb_338 = 8'h0;
  end
  if (reset) begin
    btb_339 = 8'h0;
  end
  if (reset) begin
    btb_340 = 8'h0;
  end
  if (reset) begin
    btb_341 = 8'h0;
  end
  if (reset) begin
    btb_342 = 8'h0;
  end
  if (reset) begin
    btb_343 = 8'h0;
  end
  if (reset) begin
    btb_344 = 8'h0;
  end
  if (reset) begin
    btb_345 = 8'h0;
  end
  if (reset) begin
    btb_346 = 8'h0;
  end
  if (reset) begin
    btb_347 = 8'h0;
  end
  if (reset) begin
    btb_348 = 8'h0;
  end
  if (reset) begin
    btb_349 = 8'h0;
  end
  if (reset) begin
    btb_350 = 8'h0;
  end
  if (reset) begin
    btb_351 = 8'h0;
  end
  if (reset) begin
    btb_352 = 8'h0;
  end
  if (reset) begin
    btb_353 = 8'h0;
  end
  if (reset) begin
    btb_354 = 8'h0;
  end
  if (reset) begin
    btb_355 = 8'h0;
  end
  if (reset) begin
    btb_356 = 8'h0;
  end
  if (reset) begin
    btb_357 = 8'h0;
  end
  if (reset) begin
    btb_358 = 8'h0;
  end
  if (reset) begin
    btb_359 = 8'h0;
  end
  if (reset) begin
    btb_360 = 8'h0;
  end
  if (reset) begin
    btb_361 = 8'h0;
  end
  if (reset) begin
    btb_362 = 8'h0;
  end
  if (reset) begin
    btb_363 = 8'h0;
  end
  if (reset) begin
    btb_364 = 8'h0;
  end
  if (reset) begin
    btb_365 = 8'h0;
  end
  if (reset) begin
    btb_366 = 8'h0;
  end
  if (reset) begin
    btb_367 = 8'h0;
  end
  if (reset) begin
    btb_368 = 8'h0;
  end
  if (reset) begin
    btb_369 = 8'h0;
  end
  if (reset) begin
    btb_370 = 8'h0;
  end
  if (reset) begin
    btb_371 = 8'h0;
  end
  if (reset) begin
    btb_372 = 8'h0;
  end
  if (reset) begin
    btb_373 = 8'h0;
  end
  if (reset) begin
    btb_374 = 8'h0;
  end
  if (reset) begin
    btb_375 = 8'h0;
  end
  if (reset) begin
    btb_376 = 8'h0;
  end
  if (reset) begin
    btb_377 = 8'h0;
  end
  if (reset) begin
    btb_378 = 8'h0;
  end
  if (reset) begin
    btb_379 = 8'h0;
  end
  if (reset) begin
    btb_380 = 8'h0;
  end
  if (reset) begin
    btb_381 = 8'h0;
  end
  if (reset) begin
    btb_382 = 8'h0;
  end
  if (reset) begin
    btb_383 = 8'h0;
  end
  if (reset) begin
    btb_384 = 8'h0;
  end
  if (reset) begin
    btb_385 = 8'h0;
  end
  if (reset) begin
    btb_386 = 8'h0;
  end
  if (reset) begin
    btb_387 = 8'h0;
  end
  if (reset) begin
    btb_388 = 8'h0;
  end
  if (reset) begin
    btb_389 = 8'h0;
  end
  if (reset) begin
    btb_390 = 8'h0;
  end
  if (reset) begin
    btb_391 = 8'h0;
  end
  if (reset) begin
    btb_392 = 8'h0;
  end
  if (reset) begin
    btb_393 = 8'h0;
  end
  if (reset) begin
    btb_394 = 8'h0;
  end
  if (reset) begin
    btb_395 = 8'h0;
  end
  if (reset) begin
    btb_396 = 8'h0;
  end
  if (reset) begin
    btb_397 = 8'h0;
  end
  if (reset) begin
    btb_398 = 8'h0;
  end
  if (reset) begin
    btb_399 = 8'h0;
  end
  if (reset) begin
    btb_400 = 8'h0;
  end
  if (reset) begin
    btb_401 = 8'h0;
  end
  if (reset) begin
    btb_402 = 8'h0;
  end
  if (reset) begin
    btb_403 = 8'h0;
  end
  if (reset) begin
    btb_404 = 8'h0;
  end
  if (reset) begin
    btb_405 = 8'h0;
  end
  if (reset) begin
    btb_406 = 8'h0;
  end
  if (reset) begin
    btb_407 = 8'h0;
  end
  if (reset) begin
    btb_408 = 8'h0;
  end
  if (reset) begin
    btb_409 = 8'h0;
  end
  if (reset) begin
    btb_410 = 8'h0;
  end
  if (reset) begin
    btb_411 = 8'h0;
  end
  if (reset) begin
    btb_412 = 8'h0;
  end
  if (reset) begin
    btb_413 = 8'h0;
  end
  if (reset) begin
    btb_414 = 8'h0;
  end
  if (reset) begin
    btb_415 = 8'h0;
  end
  if (reset) begin
    btb_416 = 8'h0;
  end
  if (reset) begin
    btb_417 = 8'h0;
  end
  if (reset) begin
    btb_418 = 8'h0;
  end
  if (reset) begin
    btb_419 = 8'h0;
  end
  if (reset) begin
    btb_420 = 8'h0;
  end
  if (reset) begin
    btb_421 = 8'h0;
  end
  if (reset) begin
    btb_422 = 8'h0;
  end
  if (reset) begin
    btb_423 = 8'h0;
  end
  if (reset) begin
    btb_424 = 8'h0;
  end
  if (reset) begin
    btb_425 = 8'h0;
  end
  if (reset) begin
    btb_426 = 8'h0;
  end
  if (reset) begin
    btb_427 = 8'h0;
  end
  if (reset) begin
    btb_428 = 8'h0;
  end
  if (reset) begin
    btb_429 = 8'h0;
  end
  if (reset) begin
    btb_430 = 8'h0;
  end
  if (reset) begin
    btb_431 = 8'h0;
  end
  if (reset) begin
    btb_432 = 8'h0;
  end
  if (reset) begin
    btb_433 = 8'h0;
  end
  if (reset) begin
    btb_434 = 8'h0;
  end
  if (reset) begin
    btb_435 = 8'h0;
  end
  if (reset) begin
    btb_436 = 8'h0;
  end
  if (reset) begin
    btb_437 = 8'h0;
  end
  if (reset) begin
    btb_438 = 8'h0;
  end
  if (reset) begin
    btb_439 = 8'h0;
  end
  if (reset) begin
    btb_440 = 8'h0;
  end
  if (reset) begin
    btb_441 = 8'h0;
  end
  if (reset) begin
    btb_442 = 8'h0;
  end
  if (reset) begin
    btb_443 = 8'h0;
  end
  if (reset) begin
    btb_444 = 8'h0;
  end
  if (reset) begin
    btb_445 = 8'h0;
  end
  if (reset) begin
    btb_446 = 8'h0;
  end
  if (reset) begin
    btb_447 = 8'h0;
  end
  if (reset) begin
    btb_448 = 8'h0;
  end
  if (reset) begin
    btb_449 = 8'h0;
  end
  if (reset) begin
    btb_450 = 8'h0;
  end
  if (reset) begin
    btb_451 = 8'h0;
  end
  if (reset) begin
    btb_452 = 8'h0;
  end
  if (reset) begin
    btb_453 = 8'h0;
  end
  if (reset) begin
    btb_454 = 8'h0;
  end
  if (reset) begin
    btb_455 = 8'h0;
  end
  if (reset) begin
    btb_456 = 8'h0;
  end
  if (reset) begin
    btb_457 = 8'h0;
  end
  if (reset) begin
    btb_458 = 8'h0;
  end
  if (reset) begin
    btb_459 = 8'h0;
  end
  if (reset) begin
    btb_460 = 8'h0;
  end
  if (reset) begin
    btb_461 = 8'h0;
  end
  if (reset) begin
    btb_462 = 8'h0;
  end
  if (reset) begin
    btb_463 = 8'h0;
  end
  if (reset) begin
    btb_464 = 8'h0;
  end
  if (reset) begin
    btb_465 = 8'h0;
  end
  if (reset) begin
    btb_466 = 8'h0;
  end
  if (reset) begin
    btb_467 = 8'h0;
  end
  if (reset) begin
    btb_468 = 8'h0;
  end
  if (reset) begin
    btb_469 = 8'h0;
  end
  if (reset) begin
    btb_470 = 8'h0;
  end
  if (reset) begin
    btb_471 = 8'h0;
  end
  if (reset) begin
    btb_472 = 8'h0;
  end
  if (reset) begin
    btb_473 = 8'h0;
  end
  if (reset) begin
    btb_474 = 8'h0;
  end
  if (reset) begin
    btb_475 = 8'h0;
  end
  if (reset) begin
    btb_476 = 8'h0;
  end
  if (reset) begin
    btb_477 = 8'h0;
  end
  if (reset) begin
    btb_478 = 8'h0;
  end
  if (reset) begin
    btb_479 = 8'h0;
  end
  if (reset) begin
    btb_480 = 8'h0;
  end
  if (reset) begin
    btb_481 = 8'h0;
  end
  if (reset) begin
    btb_482 = 8'h0;
  end
  if (reset) begin
    btb_483 = 8'h0;
  end
  if (reset) begin
    btb_484 = 8'h0;
  end
  if (reset) begin
    btb_485 = 8'h0;
  end
  if (reset) begin
    btb_486 = 8'h0;
  end
  if (reset) begin
    btb_487 = 8'h0;
  end
  if (reset) begin
    btb_488 = 8'h0;
  end
  if (reset) begin
    btb_489 = 8'h0;
  end
  if (reset) begin
    btb_490 = 8'h0;
  end
  if (reset) begin
    btb_491 = 8'h0;
  end
  if (reset) begin
    btb_492 = 8'h0;
  end
  if (reset) begin
    btb_493 = 8'h0;
  end
  if (reset) begin
    btb_494 = 8'h0;
  end
  if (reset) begin
    btb_495 = 8'h0;
  end
  if (reset) begin
    btb_496 = 8'h0;
  end
  if (reset) begin
    btb_497 = 8'h0;
  end
  if (reset) begin
    btb_498 = 8'h0;
  end
  if (reset) begin
    btb_499 = 8'h0;
  end
  if (reset) begin
    btb_500 = 8'h0;
  end
  if (reset) begin
    btb_501 = 8'h0;
  end
  if (reset) begin
    btb_502 = 8'h0;
  end
  if (reset) begin
    btb_503 = 8'h0;
  end
  if (reset) begin
    btb_504 = 8'h0;
  end
  if (reset) begin
    btb_505 = 8'h0;
  end
  if (reset) begin
    btb_506 = 8'h0;
  end
  if (reset) begin
    btb_507 = 8'h0;
  end
  if (reset) begin
    btb_508 = 8'h0;
  end
  if (reset) begin
    btb_509 = 8'h0;
  end
  if (reset) begin
    btb_510 = 8'h0;
  end
  if (reset) begin
    btb_511 = 8'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module data_ram_simple_two_ports_32(
  input        clock,
  input        reset,
  input        io_wea,
  input  [8:0] io_addra,
  input  [7:0] io_dina,
  input  [8:0] io_addrb,
  output [7:0] io_doutb
);
  wire  Look_up_table_read_first__clock; // @[ip_user.scala 97:23]
  wire  Look_up_table_read_first__reset; // @[ip_user.scala 97:23]
  wire [8:0] Look_up_table_read_first__io_ar_addr; // @[ip_user.scala 97:23]
  wire [8:0] Look_up_table_read_first__io_aw_addr; // @[ip_user.scala 97:23]
  wire  Look_up_table_read_first__io_write; // @[ip_user.scala 97:23]
  wire [7:0] Look_up_table_read_first__io_in; // @[ip_user.scala 97:23]
  wire [7:0] Look_up_table_read_first__io_out; // @[ip_user.scala 97:23]
  Look_up_table_read_first__32 Look_up_table_read_first_ ( // @[ip_user.scala 97:23]
    .clock(Look_up_table_read_first__clock),
    .reset(Look_up_table_read_first__reset),
    .io_ar_addr(Look_up_table_read_first__io_ar_addr),
    .io_aw_addr(Look_up_table_read_first__io_aw_addr),
    .io_write(Look_up_table_read_first__io_write),
    .io_in(Look_up_table_read_first__io_in),
    .io_out(Look_up_table_read_first__io_out)
  );
  assign io_doutb = Look_up_table_read_first__io_out; // @[ip_user.scala 102:19]
  assign Look_up_table_read_first__clock = clock;
  assign Look_up_table_read_first__reset = reset;
  assign Look_up_table_read_first__io_ar_addr = io_addra; // @[ip_user.scala 98:19]
  assign Look_up_table_read_first__io_aw_addr = io_addrb; // @[ip_user.scala 99:19]
  assign Look_up_table_read_first__io_write = io_wea; // @[ip_user.scala 101:19]
  assign Look_up_table_read_first__io_in = io_dina; // @[ip_user.scala 100:19]
endmodule
module btb_tag_with_block_ram(
  input        clock,
  input        reset,
  input        io_wen,
  input  [8:0] io_raddr,
  input  [8:0] io_waddr,
  input  [7:0] io_wdata,
  output [7:0] io_rdata
);
  wire  btb_tag_ram_0_clock; // @[BTB.scala 216:31]
  wire  btb_tag_ram_0_reset; // @[BTB.scala 216:31]
  wire  btb_tag_ram_0_io_wea; // @[BTB.scala 216:31]
  wire [8:0] btb_tag_ram_0_io_addra; // @[BTB.scala 216:31]
  wire [7:0] btb_tag_ram_0_io_dina; // @[BTB.scala 216:31]
  wire [8:0] btb_tag_ram_0_io_addrb; // @[BTB.scala 216:31]
  wire [7:0] btb_tag_ram_0_io_doutb; // @[BTB.scala 216:31]
  data_ram_simple_two_ports_32 btb_tag_ram_0 ( // @[BTB.scala 216:31]
    .clock(btb_tag_ram_0_clock),
    .reset(btb_tag_ram_0_reset),
    .io_wea(btb_tag_ram_0_io_wea),
    .io_addra(btb_tag_ram_0_io_addra),
    .io_dina(btb_tag_ram_0_io_dina),
    .io_addrb(btb_tag_ram_0_io_addrb),
    .io_doutb(btb_tag_ram_0_io_doutb)
  );
  assign io_rdata = btb_tag_ram_0_io_doutb; // @[BTB.scala 225:18]
  assign btb_tag_ram_0_clock = clock;
  assign btb_tag_ram_0_reset = reset;
  assign btb_tag_ram_0_io_wea = io_wen; // @[BTB.scala 221:27]
  assign btb_tag_ram_0_io_addra = io_waddr; // @[BTB.scala 222:28]
  assign btb_tag_ram_0_io_dina = io_wdata; // @[BTB.scala 224:27]
  assign btb_tag_ram_0_io_addrb = io_raddr; // @[BTB.scala 223:28]
endmodule
module Look_up_table_read_first__36(
  input         clock,
  input         reset,
  input  [8:0]  io_ar_addr,
  input  [8:0]  io_aw_addr,
  input         io_write,
  input  [31:0] io_in,
  output [31:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] btb_0; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_1; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_2; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_3; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_4; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_5; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_6; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_7; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_8; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_9; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_10; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_11; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_12; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_13; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_14; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_15; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_16; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_17; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_18; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_19; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_20; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_21; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_22; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_23; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_24; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_25; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_26; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_27; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_28; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_29; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_30; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_31; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_32; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_33; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_34; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_35; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_36; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_37; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_38; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_39; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_40; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_41; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_42; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_43; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_44; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_45; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_46; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_47; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_48; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_49; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_50; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_51; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_52; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_53; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_54; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_55; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_56; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_57; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_58; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_59; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_60; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_61; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_62; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_63; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_64; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_65; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_66; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_67; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_68; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_69; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_70; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_71; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_72; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_73; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_74; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_75; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_76; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_77; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_78; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_79; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_80; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_81; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_82; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_83; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_84; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_85; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_86; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_87; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_88; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_89; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_90; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_91; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_92; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_93; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_94; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_95; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_96; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_97; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_98; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_99; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_100; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_101; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_102; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_103; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_104; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_105; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_106; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_107; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_108; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_109; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_110; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_111; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_112; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_113; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_114; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_115; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_116; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_117; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_118; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_119; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_120; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_121; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_122; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_123; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_124; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_125; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_126; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_127; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_128; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_129; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_130; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_131; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_132; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_133; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_134; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_135; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_136; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_137; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_138; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_139; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_140; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_141; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_142; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_143; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_144; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_145; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_146; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_147; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_148; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_149; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_150; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_151; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_152; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_153; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_154; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_155; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_156; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_157; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_158; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_159; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_160; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_161; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_162; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_163; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_164; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_165; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_166; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_167; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_168; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_169; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_170; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_171; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_172; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_173; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_174; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_175; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_176; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_177; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_178; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_179; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_180; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_181; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_182; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_183; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_184; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_185; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_186; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_187; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_188; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_189; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_190; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_191; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_192; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_193; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_194; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_195; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_196; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_197; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_198; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_199; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_200; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_201; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_202; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_203; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_204; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_205; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_206; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_207; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_208; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_209; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_210; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_211; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_212; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_213; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_214; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_215; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_216; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_217; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_218; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_219; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_220; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_221; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_222; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_223; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_224; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_225; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_226; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_227; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_228; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_229; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_230; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_231; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_232; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_233; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_234; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_235; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_236; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_237; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_238; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_239; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_240; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_241; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_242; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_243; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_244; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_245; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_246; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_247; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_248; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_249; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_250; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_251; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_252; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_253; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_254; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_255; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_256; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_257; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_258; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_259; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_260; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_261; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_262; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_263; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_264; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_265; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_266; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_267; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_268; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_269; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_270; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_271; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_272; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_273; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_274; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_275; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_276; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_277; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_278; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_279; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_280; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_281; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_282; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_283; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_284; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_285; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_286; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_287; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_288; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_289; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_290; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_291; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_292; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_293; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_294; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_295; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_296; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_297; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_298; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_299; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_300; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_301; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_302; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_303; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_304; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_305; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_306; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_307; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_308; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_309; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_310; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_311; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_312; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_313; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_314; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_315; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_316; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_317; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_318; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_319; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_320; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_321; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_322; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_323; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_324; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_325; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_326; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_327; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_328; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_329; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_330; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_331; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_332; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_333; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_334; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_335; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_336; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_337; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_338; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_339; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_340; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_341; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_342; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_343; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_344; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_345; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_346; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_347; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_348; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_349; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_350; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_351; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_352; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_353; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_354; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_355; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_356; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_357; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_358; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_359; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_360; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_361; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_362; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_363; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_364; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_365; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_366; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_367; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_368; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_369; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_370; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_371; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_372; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_373; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_374; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_375; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_376; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_377; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_378; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_379; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_380; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_381; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_382; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_383; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_384; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_385; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_386; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_387; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_388; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_389; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_390; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_391; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_392; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_393; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_394; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_395; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_396; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_397; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_398; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_399; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_400; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_401; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_402; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_403; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_404; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_405; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_406; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_407; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_408; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_409; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_410; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_411; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_412; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_413; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_414; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_415; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_416; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_417; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_418; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_419; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_420; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_421; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_422; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_423; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_424; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_425; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_426; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_427; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_428; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_429; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_430; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_431; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_432; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_433; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_434; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_435; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_436; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_437; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_438; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_439; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_440; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_441; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_442; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_443; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_444; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_445; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_446; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_447; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_448; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_449; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_450; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_451; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_452; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_453; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_454; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_455; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_456; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_457; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_458; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_459; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_460; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_461; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_462; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_463; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_464; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_465; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_466; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_467; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_468; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_469; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_470; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_471; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_472; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_473; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_474; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_475; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_476; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_477; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_478; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_479; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_480; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_481; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_482; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_483; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_484; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_485; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_486; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_487; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_488; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_489; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_490; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_491; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_492; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_493; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_494; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_495; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_496; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_497; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_498; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_499; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_500; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_501; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_502; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_503; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_504; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_505; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_506; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_507; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_508; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_509; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_510; // @[ports_lookup_table.scala 81:22]
  reg [31:0] btb_511; // @[ports_lookup_table.scala 81:22]
  wire [31:0] _GEN_1 = 9'h1 == io_ar_addr ? btb_1 : btb_0; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_2 = 9'h2 == io_ar_addr ? btb_2 : _GEN_1; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_3 = 9'h3 == io_ar_addr ? btb_3 : _GEN_2; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_4 = 9'h4 == io_ar_addr ? btb_4 : _GEN_3; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_5 = 9'h5 == io_ar_addr ? btb_5 : _GEN_4; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_6 = 9'h6 == io_ar_addr ? btb_6 : _GEN_5; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_7 = 9'h7 == io_ar_addr ? btb_7 : _GEN_6; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_8 = 9'h8 == io_ar_addr ? btb_8 : _GEN_7; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_9 = 9'h9 == io_ar_addr ? btb_9 : _GEN_8; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_10 = 9'ha == io_ar_addr ? btb_10 : _GEN_9; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_11 = 9'hb == io_ar_addr ? btb_11 : _GEN_10; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_12 = 9'hc == io_ar_addr ? btb_12 : _GEN_11; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_13 = 9'hd == io_ar_addr ? btb_13 : _GEN_12; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_14 = 9'he == io_ar_addr ? btb_14 : _GEN_13; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_15 = 9'hf == io_ar_addr ? btb_15 : _GEN_14; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_16 = 9'h10 == io_ar_addr ? btb_16 : _GEN_15; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_17 = 9'h11 == io_ar_addr ? btb_17 : _GEN_16; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_18 = 9'h12 == io_ar_addr ? btb_18 : _GEN_17; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_19 = 9'h13 == io_ar_addr ? btb_19 : _GEN_18; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_20 = 9'h14 == io_ar_addr ? btb_20 : _GEN_19; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_21 = 9'h15 == io_ar_addr ? btb_21 : _GEN_20; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_22 = 9'h16 == io_ar_addr ? btb_22 : _GEN_21; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_23 = 9'h17 == io_ar_addr ? btb_23 : _GEN_22; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_24 = 9'h18 == io_ar_addr ? btb_24 : _GEN_23; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_25 = 9'h19 == io_ar_addr ? btb_25 : _GEN_24; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_26 = 9'h1a == io_ar_addr ? btb_26 : _GEN_25; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_27 = 9'h1b == io_ar_addr ? btb_27 : _GEN_26; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_28 = 9'h1c == io_ar_addr ? btb_28 : _GEN_27; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_29 = 9'h1d == io_ar_addr ? btb_29 : _GEN_28; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_30 = 9'h1e == io_ar_addr ? btb_30 : _GEN_29; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_31 = 9'h1f == io_ar_addr ? btb_31 : _GEN_30; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_32 = 9'h20 == io_ar_addr ? btb_32 : _GEN_31; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_33 = 9'h21 == io_ar_addr ? btb_33 : _GEN_32; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_34 = 9'h22 == io_ar_addr ? btb_34 : _GEN_33; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_35 = 9'h23 == io_ar_addr ? btb_35 : _GEN_34; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_36 = 9'h24 == io_ar_addr ? btb_36 : _GEN_35; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_37 = 9'h25 == io_ar_addr ? btb_37 : _GEN_36; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_38 = 9'h26 == io_ar_addr ? btb_38 : _GEN_37; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_39 = 9'h27 == io_ar_addr ? btb_39 : _GEN_38; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_40 = 9'h28 == io_ar_addr ? btb_40 : _GEN_39; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_41 = 9'h29 == io_ar_addr ? btb_41 : _GEN_40; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_42 = 9'h2a == io_ar_addr ? btb_42 : _GEN_41; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_43 = 9'h2b == io_ar_addr ? btb_43 : _GEN_42; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_44 = 9'h2c == io_ar_addr ? btb_44 : _GEN_43; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_45 = 9'h2d == io_ar_addr ? btb_45 : _GEN_44; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_46 = 9'h2e == io_ar_addr ? btb_46 : _GEN_45; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_47 = 9'h2f == io_ar_addr ? btb_47 : _GEN_46; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_48 = 9'h30 == io_ar_addr ? btb_48 : _GEN_47; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_49 = 9'h31 == io_ar_addr ? btb_49 : _GEN_48; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_50 = 9'h32 == io_ar_addr ? btb_50 : _GEN_49; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_51 = 9'h33 == io_ar_addr ? btb_51 : _GEN_50; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_52 = 9'h34 == io_ar_addr ? btb_52 : _GEN_51; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_53 = 9'h35 == io_ar_addr ? btb_53 : _GEN_52; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_54 = 9'h36 == io_ar_addr ? btb_54 : _GEN_53; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_55 = 9'h37 == io_ar_addr ? btb_55 : _GEN_54; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_56 = 9'h38 == io_ar_addr ? btb_56 : _GEN_55; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_57 = 9'h39 == io_ar_addr ? btb_57 : _GEN_56; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_58 = 9'h3a == io_ar_addr ? btb_58 : _GEN_57; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_59 = 9'h3b == io_ar_addr ? btb_59 : _GEN_58; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_60 = 9'h3c == io_ar_addr ? btb_60 : _GEN_59; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_61 = 9'h3d == io_ar_addr ? btb_61 : _GEN_60; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_62 = 9'h3e == io_ar_addr ? btb_62 : _GEN_61; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_63 = 9'h3f == io_ar_addr ? btb_63 : _GEN_62; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_64 = 9'h40 == io_ar_addr ? btb_64 : _GEN_63; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_65 = 9'h41 == io_ar_addr ? btb_65 : _GEN_64; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_66 = 9'h42 == io_ar_addr ? btb_66 : _GEN_65; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_67 = 9'h43 == io_ar_addr ? btb_67 : _GEN_66; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_68 = 9'h44 == io_ar_addr ? btb_68 : _GEN_67; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_69 = 9'h45 == io_ar_addr ? btb_69 : _GEN_68; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_70 = 9'h46 == io_ar_addr ? btb_70 : _GEN_69; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_71 = 9'h47 == io_ar_addr ? btb_71 : _GEN_70; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_72 = 9'h48 == io_ar_addr ? btb_72 : _GEN_71; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_73 = 9'h49 == io_ar_addr ? btb_73 : _GEN_72; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_74 = 9'h4a == io_ar_addr ? btb_74 : _GEN_73; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_75 = 9'h4b == io_ar_addr ? btb_75 : _GEN_74; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_76 = 9'h4c == io_ar_addr ? btb_76 : _GEN_75; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_77 = 9'h4d == io_ar_addr ? btb_77 : _GEN_76; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_78 = 9'h4e == io_ar_addr ? btb_78 : _GEN_77; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_79 = 9'h4f == io_ar_addr ? btb_79 : _GEN_78; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_80 = 9'h50 == io_ar_addr ? btb_80 : _GEN_79; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_81 = 9'h51 == io_ar_addr ? btb_81 : _GEN_80; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_82 = 9'h52 == io_ar_addr ? btb_82 : _GEN_81; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_83 = 9'h53 == io_ar_addr ? btb_83 : _GEN_82; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_84 = 9'h54 == io_ar_addr ? btb_84 : _GEN_83; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_85 = 9'h55 == io_ar_addr ? btb_85 : _GEN_84; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_86 = 9'h56 == io_ar_addr ? btb_86 : _GEN_85; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_87 = 9'h57 == io_ar_addr ? btb_87 : _GEN_86; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_88 = 9'h58 == io_ar_addr ? btb_88 : _GEN_87; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_89 = 9'h59 == io_ar_addr ? btb_89 : _GEN_88; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_90 = 9'h5a == io_ar_addr ? btb_90 : _GEN_89; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_91 = 9'h5b == io_ar_addr ? btb_91 : _GEN_90; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_92 = 9'h5c == io_ar_addr ? btb_92 : _GEN_91; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_93 = 9'h5d == io_ar_addr ? btb_93 : _GEN_92; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_94 = 9'h5e == io_ar_addr ? btb_94 : _GEN_93; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_95 = 9'h5f == io_ar_addr ? btb_95 : _GEN_94; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_96 = 9'h60 == io_ar_addr ? btb_96 : _GEN_95; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_97 = 9'h61 == io_ar_addr ? btb_97 : _GEN_96; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_98 = 9'h62 == io_ar_addr ? btb_98 : _GEN_97; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_99 = 9'h63 == io_ar_addr ? btb_99 : _GEN_98; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_100 = 9'h64 == io_ar_addr ? btb_100 : _GEN_99; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_101 = 9'h65 == io_ar_addr ? btb_101 : _GEN_100; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_102 = 9'h66 == io_ar_addr ? btb_102 : _GEN_101; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_103 = 9'h67 == io_ar_addr ? btb_103 : _GEN_102; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_104 = 9'h68 == io_ar_addr ? btb_104 : _GEN_103; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_105 = 9'h69 == io_ar_addr ? btb_105 : _GEN_104; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_106 = 9'h6a == io_ar_addr ? btb_106 : _GEN_105; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_107 = 9'h6b == io_ar_addr ? btb_107 : _GEN_106; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_108 = 9'h6c == io_ar_addr ? btb_108 : _GEN_107; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_109 = 9'h6d == io_ar_addr ? btb_109 : _GEN_108; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_110 = 9'h6e == io_ar_addr ? btb_110 : _GEN_109; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_111 = 9'h6f == io_ar_addr ? btb_111 : _GEN_110; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_112 = 9'h70 == io_ar_addr ? btb_112 : _GEN_111; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_113 = 9'h71 == io_ar_addr ? btb_113 : _GEN_112; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_114 = 9'h72 == io_ar_addr ? btb_114 : _GEN_113; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_115 = 9'h73 == io_ar_addr ? btb_115 : _GEN_114; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_116 = 9'h74 == io_ar_addr ? btb_116 : _GEN_115; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_117 = 9'h75 == io_ar_addr ? btb_117 : _GEN_116; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_118 = 9'h76 == io_ar_addr ? btb_118 : _GEN_117; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_119 = 9'h77 == io_ar_addr ? btb_119 : _GEN_118; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_120 = 9'h78 == io_ar_addr ? btb_120 : _GEN_119; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_121 = 9'h79 == io_ar_addr ? btb_121 : _GEN_120; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_122 = 9'h7a == io_ar_addr ? btb_122 : _GEN_121; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_123 = 9'h7b == io_ar_addr ? btb_123 : _GEN_122; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_124 = 9'h7c == io_ar_addr ? btb_124 : _GEN_123; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_125 = 9'h7d == io_ar_addr ? btb_125 : _GEN_124; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_126 = 9'h7e == io_ar_addr ? btb_126 : _GEN_125; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_127 = 9'h7f == io_ar_addr ? btb_127 : _GEN_126; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_128 = 9'h80 == io_ar_addr ? btb_128 : _GEN_127; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_129 = 9'h81 == io_ar_addr ? btb_129 : _GEN_128; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_130 = 9'h82 == io_ar_addr ? btb_130 : _GEN_129; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_131 = 9'h83 == io_ar_addr ? btb_131 : _GEN_130; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_132 = 9'h84 == io_ar_addr ? btb_132 : _GEN_131; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_133 = 9'h85 == io_ar_addr ? btb_133 : _GEN_132; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_134 = 9'h86 == io_ar_addr ? btb_134 : _GEN_133; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_135 = 9'h87 == io_ar_addr ? btb_135 : _GEN_134; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_136 = 9'h88 == io_ar_addr ? btb_136 : _GEN_135; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_137 = 9'h89 == io_ar_addr ? btb_137 : _GEN_136; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_138 = 9'h8a == io_ar_addr ? btb_138 : _GEN_137; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_139 = 9'h8b == io_ar_addr ? btb_139 : _GEN_138; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_140 = 9'h8c == io_ar_addr ? btb_140 : _GEN_139; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_141 = 9'h8d == io_ar_addr ? btb_141 : _GEN_140; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_142 = 9'h8e == io_ar_addr ? btb_142 : _GEN_141; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_143 = 9'h8f == io_ar_addr ? btb_143 : _GEN_142; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_144 = 9'h90 == io_ar_addr ? btb_144 : _GEN_143; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_145 = 9'h91 == io_ar_addr ? btb_145 : _GEN_144; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_146 = 9'h92 == io_ar_addr ? btb_146 : _GEN_145; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_147 = 9'h93 == io_ar_addr ? btb_147 : _GEN_146; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_148 = 9'h94 == io_ar_addr ? btb_148 : _GEN_147; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_149 = 9'h95 == io_ar_addr ? btb_149 : _GEN_148; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_150 = 9'h96 == io_ar_addr ? btb_150 : _GEN_149; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_151 = 9'h97 == io_ar_addr ? btb_151 : _GEN_150; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_152 = 9'h98 == io_ar_addr ? btb_152 : _GEN_151; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_153 = 9'h99 == io_ar_addr ? btb_153 : _GEN_152; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_154 = 9'h9a == io_ar_addr ? btb_154 : _GEN_153; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_155 = 9'h9b == io_ar_addr ? btb_155 : _GEN_154; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_156 = 9'h9c == io_ar_addr ? btb_156 : _GEN_155; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_157 = 9'h9d == io_ar_addr ? btb_157 : _GEN_156; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_158 = 9'h9e == io_ar_addr ? btb_158 : _GEN_157; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_159 = 9'h9f == io_ar_addr ? btb_159 : _GEN_158; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_160 = 9'ha0 == io_ar_addr ? btb_160 : _GEN_159; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_161 = 9'ha1 == io_ar_addr ? btb_161 : _GEN_160; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_162 = 9'ha2 == io_ar_addr ? btb_162 : _GEN_161; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_163 = 9'ha3 == io_ar_addr ? btb_163 : _GEN_162; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_164 = 9'ha4 == io_ar_addr ? btb_164 : _GEN_163; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_165 = 9'ha5 == io_ar_addr ? btb_165 : _GEN_164; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_166 = 9'ha6 == io_ar_addr ? btb_166 : _GEN_165; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_167 = 9'ha7 == io_ar_addr ? btb_167 : _GEN_166; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_168 = 9'ha8 == io_ar_addr ? btb_168 : _GEN_167; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_169 = 9'ha9 == io_ar_addr ? btb_169 : _GEN_168; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_170 = 9'haa == io_ar_addr ? btb_170 : _GEN_169; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_171 = 9'hab == io_ar_addr ? btb_171 : _GEN_170; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_172 = 9'hac == io_ar_addr ? btb_172 : _GEN_171; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_173 = 9'had == io_ar_addr ? btb_173 : _GEN_172; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_174 = 9'hae == io_ar_addr ? btb_174 : _GEN_173; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_175 = 9'haf == io_ar_addr ? btb_175 : _GEN_174; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_176 = 9'hb0 == io_ar_addr ? btb_176 : _GEN_175; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_177 = 9'hb1 == io_ar_addr ? btb_177 : _GEN_176; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_178 = 9'hb2 == io_ar_addr ? btb_178 : _GEN_177; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_179 = 9'hb3 == io_ar_addr ? btb_179 : _GEN_178; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_180 = 9'hb4 == io_ar_addr ? btb_180 : _GEN_179; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_181 = 9'hb5 == io_ar_addr ? btb_181 : _GEN_180; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_182 = 9'hb6 == io_ar_addr ? btb_182 : _GEN_181; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_183 = 9'hb7 == io_ar_addr ? btb_183 : _GEN_182; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_184 = 9'hb8 == io_ar_addr ? btb_184 : _GEN_183; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_185 = 9'hb9 == io_ar_addr ? btb_185 : _GEN_184; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_186 = 9'hba == io_ar_addr ? btb_186 : _GEN_185; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_187 = 9'hbb == io_ar_addr ? btb_187 : _GEN_186; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_188 = 9'hbc == io_ar_addr ? btb_188 : _GEN_187; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_189 = 9'hbd == io_ar_addr ? btb_189 : _GEN_188; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_190 = 9'hbe == io_ar_addr ? btb_190 : _GEN_189; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_191 = 9'hbf == io_ar_addr ? btb_191 : _GEN_190; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_192 = 9'hc0 == io_ar_addr ? btb_192 : _GEN_191; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_193 = 9'hc1 == io_ar_addr ? btb_193 : _GEN_192; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_194 = 9'hc2 == io_ar_addr ? btb_194 : _GEN_193; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_195 = 9'hc3 == io_ar_addr ? btb_195 : _GEN_194; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_196 = 9'hc4 == io_ar_addr ? btb_196 : _GEN_195; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_197 = 9'hc5 == io_ar_addr ? btb_197 : _GEN_196; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_198 = 9'hc6 == io_ar_addr ? btb_198 : _GEN_197; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_199 = 9'hc7 == io_ar_addr ? btb_199 : _GEN_198; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_200 = 9'hc8 == io_ar_addr ? btb_200 : _GEN_199; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_201 = 9'hc9 == io_ar_addr ? btb_201 : _GEN_200; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_202 = 9'hca == io_ar_addr ? btb_202 : _GEN_201; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_203 = 9'hcb == io_ar_addr ? btb_203 : _GEN_202; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_204 = 9'hcc == io_ar_addr ? btb_204 : _GEN_203; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_205 = 9'hcd == io_ar_addr ? btb_205 : _GEN_204; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_206 = 9'hce == io_ar_addr ? btb_206 : _GEN_205; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_207 = 9'hcf == io_ar_addr ? btb_207 : _GEN_206; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_208 = 9'hd0 == io_ar_addr ? btb_208 : _GEN_207; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_209 = 9'hd1 == io_ar_addr ? btb_209 : _GEN_208; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_210 = 9'hd2 == io_ar_addr ? btb_210 : _GEN_209; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_211 = 9'hd3 == io_ar_addr ? btb_211 : _GEN_210; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_212 = 9'hd4 == io_ar_addr ? btb_212 : _GEN_211; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_213 = 9'hd5 == io_ar_addr ? btb_213 : _GEN_212; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_214 = 9'hd6 == io_ar_addr ? btb_214 : _GEN_213; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_215 = 9'hd7 == io_ar_addr ? btb_215 : _GEN_214; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_216 = 9'hd8 == io_ar_addr ? btb_216 : _GEN_215; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_217 = 9'hd9 == io_ar_addr ? btb_217 : _GEN_216; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_218 = 9'hda == io_ar_addr ? btb_218 : _GEN_217; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_219 = 9'hdb == io_ar_addr ? btb_219 : _GEN_218; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_220 = 9'hdc == io_ar_addr ? btb_220 : _GEN_219; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_221 = 9'hdd == io_ar_addr ? btb_221 : _GEN_220; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_222 = 9'hde == io_ar_addr ? btb_222 : _GEN_221; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_223 = 9'hdf == io_ar_addr ? btb_223 : _GEN_222; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_224 = 9'he0 == io_ar_addr ? btb_224 : _GEN_223; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_225 = 9'he1 == io_ar_addr ? btb_225 : _GEN_224; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_226 = 9'he2 == io_ar_addr ? btb_226 : _GEN_225; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_227 = 9'he3 == io_ar_addr ? btb_227 : _GEN_226; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_228 = 9'he4 == io_ar_addr ? btb_228 : _GEN_227; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_229 = 9'he5 == io_ar_addr ? btb_229 : _GEN_228; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_230 = 9'he6 == io_ar_addr ? btb_230 : _GEN_229; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_231 = 9'he7 == io_ar_addr ? btb_231 : _GEN_230; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_232 = 9'he8 == io_ar_addr ? btb_232 : _GEN_231; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_233 = 9'he9 == io_ar_addr ? btb_233 : _GEN_232; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_234 = 9'hea == io_ar_addr ? btb_234 : _GEN_233; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_235 = 9'heb == io_ar_addr ? btb_235 : _GEN_234; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_236 = 9'hec == io_ar_addr ? btb_236 : _GEN_235; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_237 = 9'hed == io_ar_addr ? btb_237 : _GEN_236; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_238 = 9'hee == io_ar_addr ? btb_238 : _GEN_237; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_239 = 9'hef == io_ar_addr ? btb_239 : _GEN_238; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_240 = 9'hf0 == io_ar_addr ? btb_240 : _GEN_239; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_241 = 9'hf1 == io_ar_addr ? btb_241 : _GEN_240; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_242 = 9'hf2 == io_ar_addr ? btb_242 : _GEN_241; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_243 = 9'hf3 == io_ar_addr ? btb_243 : _GEN_242; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_244 = 9'hf4 == io_ar_addr ? btb_244 : _GEN_243; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_245 = 9'hf5 == io_ar_addr ? btb_245 : _GEN_244; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_246 = 9'hf6 == io_ar_addr ? btb_246 : _GEN_245; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_247 = 9'hf7 == io_ar_addr ? btb_247 : _GEN_246; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_248 = 9'hf8 == io_ar_addr ? btb_248 : _GEN_247; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_249 = 9'hf9 == io_ar_addr ? btb_249 : _GEN_248; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_250 = 9'hfa == io_ar_addr ? btb_250 : _GEN_249; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_251 = 9'hfb == io_ar_addr ? btb_251 : _GEN_250; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_252 = 9'hfc == io_ar_addr ? btb_252 : _GEN_251; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_253 = 9'hfd == io_ar_addr ? btb_253 : _GEN_252; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_254 = 9'hfe == io_ar_addr ? btb_254 : _GEN_253; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_255 = 9'hff == io_ar_addr ? btb_255 : _GEN_254; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_256 = 9'h100 == io_ar_addr ? btb_256 : _GEN_255; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_257 = 9'h101 == io_ar_addr ? btb_257 : _GEN_256; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_258 = 9'h102 == io_ar_addr ? btb_258 : _GEN_257; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_259 = 9'h103 == io_ar_addr ? btb_259 : _GEN_258; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_260 = 9'h104 == io_ar_addr ? btb_260 : _GEN_259; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_261 = 9'h105 == io_ar_addr ? btb_261 : _GEN_260; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_262 = 9'h106 == io_ar_addr ? btb_262 : _GEN_261; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_263 = 9'h107 == io_ar_addr ? btb_263 : _GEN_262; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_264 = 9'h108 == io_ar_addr ? btb_264 : _GEN_263; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_265 = 9'h109 == io_ar_addr ? btb_265 : _GEN_264; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_266 = 9'h10a == io_ar_addr ? btb_266 : _GEN_265; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_267 = 9'h10b == io_ar_addr ? btb_267 : _GEN_266; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_268 = 9'h10c == io_ar_addr ? btb_268 : _GEN_267; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_269 = 9'h10d == io_ar_addr ? btb_269 : _GEN_268; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_270 = 9'h10e == io_ar_addr ? btb_270 : _GEN_269; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_271 = 9'h10f == io_ar_addr ? btb_271 : _GEN_270; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_272 = 9'h110 == io_ar_addr ? btb_272 : _GEN_271; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_273 = 9'h111 == io_ar_addr ? btb_273 : _GEN_272; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_274 = 9'h112 == io_ar_addr ? btb_274 : _GEN_273; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_275 = 9'h113 == io_ar_addr ? btb_275 : _GEN_274; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_276 = 9'h114 == io_ar_addr ? btb_276 : _GEN_275; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_277 = 9'h115 == io_ar_addr ? btb_277 : _GEN_276; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_278 = 9'h116 == io_ar_addr ? btb_278 : _GEN_277; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_279 = 9'h117 == io_ar_addr ? btb_279 : _GEN_278; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_280 = 9'h118 == io_ar_addr ? btb_280 : _GEN_279; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_281 = 9'h119 == io_ar_addr ? btb_281 : _GEN_280; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_282 = 9'h11a == io_ar_addr ? btb_282 : _GEN_281; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_283 = 9'h11b == io_ar_addr ? btb_283 : _GEN_282; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_284 = 9'h11c == io_ar_addr ? btb_284 : _GEN_283; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_285 = 9'h11d == io_ar_addr ? btb_285 : _GEN_284; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_286 = 9'h11e == io_ar_addr ? btb_286 : _GEN_285; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_287 = 9'h11f == io_ar_addr ? btb_287 : _GEN_286; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_288 = 9'h120 == io_ar_addr ? btb_288 : _GEN_287; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_289 = 9'h121 == io_ar_addr ? btb_289 : _GEN_288; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_290 = 9'h122 == io_ar_addr ? btb_290 : _GEN_289; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_291 = 9'h123 == io_ar_addr ? btb_291 : _GEN_290; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_292 = 9'h124 == io_ar_addr ? btb_292 : _GEN_291; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_293 = 9'h125 == io_ar_addr ? btb_293 : _GEN_292; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_294 = 9'h126 == io_ar_addr ? btb_294 : _GEN_293; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_295 = 9'h127 == io_ar_addr ? btb_295 : _GEN_294; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_296 = 9'h128 == io_ar_addr ? btb_296 : _GEN_295; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_297 = 9'h129 == io_ar_addr ? btb_297 : _GEN_296; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_298 = 9'h12a == io_ar_addr ? btb_298 : _GEN_297; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_299 = 9'h12b == io_ar_addr ? btb_299 : _GEN_298; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_300 = 9'h12c == io_ar_addr ? btb_300 : _GEN_299; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_301 = 9'h12d == io_ar_addr ? btb_301 : _GEN_300; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_302 = 9'h12e == io_ar_addr ? btb_302 : _GEN_301; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_303 = 9'h12f == io_ar_addr ? btb_303 : _GEN_302; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_304 = 9'h130 == io_ar_addr ? btb_304 : _GEN_303; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_305 = 9'h131 == io_ar_addr ? btb_305 : _GEN_304; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_306 = 9'h132 == io_ar_addr ? btb_306 : _GEN_305; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_307 = 9'h133 == io_ar_addr ? btb_307 : _GEN_306; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_308 = 9'h134 == io_ar_addr ? btb_308 : _GEN_307; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_309 = 9'h135 == io_ar_addr ? btb_309 : _GEN_308; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_310 = 9'h136 == io_ar_addr ? btb_310 : _GEN_309; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_311 = 9'h137 == io_ar_addr ? btb_311 : _GEN_310; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_312 = 9'h138 == io_ar_addr ? btb_312 : _GEN_311; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_313 = 9'h139 == io_ar_addr ? btb_313 : _GEN_312; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_314 = 9'h13a == io_ar_addr ? btb_314 : _GEN_313; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_315 = 9'h13b == io_ar_addr ? btb_315 : _GEN_314; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_316 = 9'h13c == io_ar_addr ? btb_316 : _GEN_315; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_317 = 9'h13d == io_ar_addr ? btb_317 : _GEN_316; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_318 = 9'h13e == io_ar_addr ? btb_318 : _GEN_317; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_319 = 9'h13f == io_ar_addr ? btb_319 : _GEN_318; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_320 = 9'h140 == io_ar_addr ? btb_320 : _GEN_319; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_321 = 9'h141 == io_ar_addr ? btb_321 : _GEN_320; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_322 = 9'h142 == io_ar_addr ? btb_322 : _GEN_321; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_323 = 9'h143 == io_ar_addr ? btb_323 : _GEN_322; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_324 = 9'h144 == io_ar_addr ? btb_324 : _GEN_323; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_325 = 9'h145 == io_ar_addr ? btb_325 : _GEN_324; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_326 = 9'h146 == io_ar_addr ? btb_326 : _GEN_325; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_327 = 9'h147 == io_ar_addr ? btb_327 : _GEN_326; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_328 = 9'h148 == io_ar_addr ? btb_328 : _GEN_327; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_329 = 9'h149 == io_ar_addr ? btb_329 : _GEN_328; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_330 = 9'h14a == io_ar_addr ? btb_330 : _GEN_329; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_331 = 9'h14b == io_ar_addr ? btb_331 : _GEN_330; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_332 = 9'h14c == io_ar_addr ? btb_332 : _GEN_331; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_333 = 9'h14d == io_ar_addr ? btb_333 : _GEN_332; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_334 = 9'h14e == io_ar_addr ? btb_334 : _GEN_333; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_335 = 9'h14f == io_ar_addr ? btb_335 : _GEN_334; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_336 = 9'h150 == io_ar_addr ? btb_336 : _GEN_335; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_337 = 9'h151 == io_ar_addr ? btb_337 : _GEN_336; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_338 = 9'h152 == io_ar_addr ? btb_338 : _GEN_337; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_339 = 9'h153 == io_ar_addr ? btb_339 : _GEN_338; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_340 = 9'h154 == io_ar_addr ? btb_340 : _GEN_339; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_341 = 9'h155 == io_ar_addr ? btb_341 : _GEN_340; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_342 = 9'h156 == io_ar_addr ? btb_342 : _GEN_341; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_343 = 9'h157 == io_ar_addr ? btb_343 : _GEN_342; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_344 = 9'h158 == io_ar_addr ? btb_344 : _GEN_343; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_345 = 9'h159 == io_ar_addr ? btb_345 : _GEN_344; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_346 = 9'h15a == io_ar_addr ? btb_346 : _GEN_345; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_347 = 9'h15b == io_ar_addr ? btb_347 : _GEN_346; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_348 = 9'h15c == io_ar_addr ? btb_348 : _GEN_347; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_349 = 9'h15d == io_ar_addr ? btb_349 : _GEN_348; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_350 = 9'h15e == io_ar_addr ? btb_350 : _GEN_349; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_351 = 9'h15f == io_ar_addr ? btb_351 : _GEN_350; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_352 = 9'h160 == io_ar_addr ? btb_352 : _GEN_351; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_353 = 9'h161 == io_ar_addr ? btb_353 : _GEN_352; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_354 = 9'h162 == io_ar_addr ? btb_354 : _GEN_353; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_355 = 9'h163 == io_ar_addr ? btb_355 : _GEN_354; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_356 = 9'h164 == io_ar_addr ? btb_356 : _GEN_355; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_357 = 9'h165 == io_ar_addr ? btb_357 : _GEN_356; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_358 = 9'h166 == io_ar_addr ? btb_358 : _GEN_357; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_359 = 9'h167 == io_ar_addr ? btb_359 : _GEN_358; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_360 = 9'h168 == io_ar_addr ? btb_360 : _GEN_359; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_361 = 9'h169 == io_ar_addr ? btb_361 : _GEN_360; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_362 = 9'h16a == io_ar_addr ? btb_362 : _GEN_361; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_363 = 9'h16b == io_ar_addr ? btb_363 : _GEN_362; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_364 = 9'h16c == io_ar_addr ? btb_364 : _GEN_363; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_365 = 9'h16d == io_ar_addr ? btb_365 : _GEN_364; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_366 = 9'h16e == io_ar_addr ? btb_366 : _GEN_365; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_367 = 9'h16f == io_ar_addr ? btb_367 : _GEN_366; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_368 = 9'h170 == io_ar_addr ? btb_368 : _GEN_367; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_369 = 9'h171 == io_ar_addr ? btb_369 : _GEN_368; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_370 = 9'h172 == io_ar_addr ? btb_370 : _GEN_369; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_371 = 9'h173 == io_ar_addr ? btb_371 : _GEN_370; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_372 = 9'h174 == io_ar_addr ? btb_372 : _GEN_371; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_373 = 9'h175 == io_ar_addr ? btb_373 : _GEN_372; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_374 = 9'h176 == io_ar_addr ? btb_374 : _GEN_373; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_375 = 9'h177 == io_ar_addr ? btb_375 : _GEN_374; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_376 = 9'h178 == io_ar_addr ? btb_376 : _GEN_375; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_377 = 9'h179 == io_ar_addr ? btb_377 : _GEN_376; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_378 = 9'h17a == io_ar_addr ? btb_378 : _GEN_377; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_379 = 9'h17b == io_ar_addr ? btb_379 : _GEN_378; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_380 = 9'h17c == io_ar_addr ? btb_380 : _GEN_379; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_381 = 9'h17d == io_ar_addr ? btb_381 : _GEN_380; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_382 = 9'h17e == io_ar_addr ? btb_382 : _GEN_381; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_383 = 9'h17f == io_ar_addr ? btb_383 : _GEN_382; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_384 = 9'h180 == io_ar_addr ? btb_384 : _GEN_383; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_385 = 9'h181 == io_ar_addr ? btb_385 : _GEN_384; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_386 = 9'h182 == io_ar_addr ? btb_386 : _GEN_385; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_387 = 9'h183 == io_ar_addr ? btb_387 : _GEN_386; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_388 = 9'h184 == io_ar_addr ? btb_388 : _GEN_387; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_389 = 9'h185 == io_ar_addr ? btb_389 : _GEN_388; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_390 = 9'h186 == io_ar_addr ? btb_390 : _GEN_389; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_391 = 9'h187 == io_ar_addr ? btb_391 : _GEN_390; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_392 = 9'h188 == io_ar_addr ? btb_392 : _GEN_391; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_393 = 9'h189 == io_ar_addr ? btb_393 : _GEN_392; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_394 = 9'h18a == io_ar_addr ? btb_394 : _GEN_393; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_395 = 9'h18b == io_ar_addr ? btb_395 : _GEN_394; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_396 = 9'h18c == io_ar_addr ? btb_396 : _GEN_395; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_397 = 9'h18d == io_ar_addr ? btb_397 : _GEN_396; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_398 = 9'h18e == io_ar_addr ? btb_398 : _GEN_397; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_399 = 9'h18f == io_ar_addr ? btb_399 : _GEN_398; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_400 = 9'h190 == io_ar_addr ? btb_400 : _GEN_399; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_401 = 9'h191 == io_ar_addr ? btb_401 : _GEN_400; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_402 = 9'h192 == io_ar_addr ? btb_402 : _GEN_401; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_403 = 9'h193 == io_ar_addr ? btb_403 : _GEN_402; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_404 = 9'h194 == io_ar_addr ? btb_404 : _GEN_403; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_405 = 9'h195 == io_ar_addr ? btb_405 : _GEN_404; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_406 = 9'h196 == io_ar_addr ? btb_406 : _GEN_405; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_407 = 9'h197 == io_ar_addr ? btb_407 : _GEN_406; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_408 = 9'h198 == io_ar_addr ? btb_408 : _GEN_407; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_409 = 9'h199 == io_ar_addr ? btb_409 : _GEN_408; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_410 = 9'h19a == io_ar_addr ? btb_410 : _GEN_409; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_411 = 9'h19b == io_ar_addr ? btb_411 : _GEN_410; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_412 = 9'h19c == io_ar_addr ? btb_412 : _GEN_411; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_413 = 9'h19d == io_ar_addr ? btb_413 : _GEN_412; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_414 = 9'h19e == io_ar_addr ? btb_414 : _GEN_413; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_415 = 9'h19f == io_ar_addr ? btb_415 : _GEN_414; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_416 = 9'h1a0 == io_ar_addr ? btb_416 : _GEN_415; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_417 = 9'h1a1 == io_ar_addr ? btb_417 : _GEN_416; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_418 = 9'h1a2 == io_ar_addr ? btb_418 : _GEN_417; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_419 = 9'h1a3 == io_ar_addr ? btb_419 : _GEN_418; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_420 = 9'h1a4 == io_ar_addr ? btb_420 : _GEN_419; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_421 = 9'h1a5 == io_ar_addr ? btb_421 : _GEN_420; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_422 = 9'h1a6 == io_ar_addr ? btb_422 : _GEN_421; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_423 = 9'h1a7 == io_ar_addr ? btb_423 : _GEN_422; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_424 = 9'h1a8 == io_ar_addr ? btb_424 : _GEN_423; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_425 = 9'h1a9 == io_ar_addr ? btb_425 : _GEN_424; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_426 = 9'h1aa == io_ar_addr ? btb_426 : _GEN_425; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_427 = 9'h1ab == io_ar_addr ? btb_427 : _GEN_426; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_428 = 9'h1ac == io_ar_addr ? btb_428 : _GEN_427; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_429 = 9'h1ad == io_ar_addr ? btb_429 : _GEN_428; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_430 = 9'h1ae == io_ar_addr ? btb_430 : _GEN_429; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_431 = 9'h1af == io_ar_addr ? btb_431 : _GEN_430; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_432 = 9'h1b0 == io_ar_addr ? btb_432 : _GEN_431; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_433 = 9'h1b1 == io_ar_addr ? btb_433 : _GEN_432; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_434 = 9'h1b2 == io_ar_addr ? btb_434 : _GEN_433; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_435 = 9'h1b3 == io_ar_addr ? btb_435 : _GEN_434; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_436 = 9'h1b4 == io_ar_addr ? btb_436 : _GEN_435; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_437 = 9'h1b5 == io_ar_addr ? btb_437 : _GEN_436; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_438 = 9'h1b6 == io_ar_addr ? btb_438 : _GEN_437; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_439 = 9'h1b7 == io_ar_addr ? btb_439 : _GEN_438; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_440 = 9'h1b8 == io_ar_addr ? btb_440 : _GEN_439; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_441 = 9'h1b9 == io_ar_addr ? btb_441 : _GEN_440; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_442 = 9'h1ba == io_ar_addr ? btb_442 : _GEN_441; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_443 = 9'h1bb == io_ar_addr ? btb_443 : _GEN_442; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_444 = 9'h1bc == io_ar_addr ? btb_444 : _GEN_443; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_445 = 9'h1bd == io_ar_addr ? btb_445 : _GEN_444; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_446 = 9'h1be == io_ar_addr ? btb_446 : _GEN_445; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_447 = 9'h1bf == io_ar_addr ? btb_447 : _GEN_446; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_448 = 9'h1c0 == io_ar_addr ? btb_448 : _GEN_447; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_449 = 9'h1c1 == io_ar_addr ? btb_449 : _GEN_448; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_450 = 9'h1c2 == io_ar_addr ? btb_450 : _GEN_449; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_451 = 9'h1c3 == io_ar_addr ? btb_451 : _GEN_450; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_452 = 9'h1c4 == io_ar_addr ? btb_452 : _GEN_451; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_453 = 9'h1c5 == io_ar_addr ? btb_453 : _GEN_452; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_454 = 9'h1c6 == io_ar_addr ? btb_454 : _GEN_453; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_455 = 9'h1c7 == io_ar_addr ? btb_455 : _GEN_454; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_456 = 9'h1c8 == io_ar_addr ? btb_456 : _GEN_455; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_457 = 9'h1c9 == io_ar_addr ? btb_457 : _GEN_456; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_458 = 9'h1ca == io_ar_addr ? btb_458 : _GEN_457; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_459 = 9'h1cb == io_ar_addr ? btb_459 : _GEN_458; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_460 = 9'h1cc == io_ar_addr ? btb_460 : _GEN_459; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_461 = 9'h1cd == io_ar_addr ? btb_461 : _GEN_460; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_462 = 9'h1ce == io_ar_addr ? btb_462 : _GEN_461; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_463 = 9'h1cf == io_ar_addr ? btb_463 : _GEN_462; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_464 = 9'h1d0 == io_ar_addr ? btb_464 : _GEN_463; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_465 = 9'h1d1 == io_ar_addr ? btb_465 : _GEN_464; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_466 = 9'h1d2 == io_ar_addr ? btb_466 : _GEN_465; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_467 = 9'h1d3 == io_ar_addr ? btb_467 : _GEN_466; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_468 = 9'h1d4 == io_ar_addr ? btb_468 : _GEN_467; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_469 = 9'h1d5 == io_ar_addr ? btb_469 : _GEN_468; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_470 = 9'h1d6 == io_ar_addr ? btb_470 : _GEN_469; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_471 = 9'h1d7 == io_ar_addr ? btb_471 : _GEN_470; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_472 = 9'h1d8 == io_ar_addr ? btb_472 : _GEN_471; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_473 = 9'h1d9 == io_ar_addr ? btb_473 : _GEN_472; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_474 = 9'h1da == io_ar_addr ? btb_474 : _GEN_473; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_475 = 9'h1db == io_ar_addr ? btb_475 : _GEN_474; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_476 = 9'h1dc == io_ar_addr ? btb_476 : _GEN_475; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_477 = 9'h1dd == io_ar_addr ? btb_477 : _GEN_476; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_478 = 9'h1de == io_ar_addr ? btb_478 : _GEN_477; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_479 = 9'h1df == io_ar_addr ? btb_479 : _GEN_478; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_480 = 9'h1e0 == io_ar_addr ? btb_480 : _GEN_479; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_481 = 9'h1e1 == io_ar_addr ? btb_481 : _GEN_480; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_482 = 9'h1e2 == io_ar_addr ? btb_482 : _GEN_481; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_483 = 9'h1e3 == io_ar_addr ? btb_483 : _GEN_482; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_484 = 9'h1e4 == io_ar_addr ? btb_484 : _GEN_483; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_485 = 9'h1e5 == io_ar_addr ? btb_485 : _GEN_484; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_486 = 9'h1e6 == io_ar_addr ? btb_486 : _GEN_485; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_487 = 9'h1e7 == io_ar_addr ? btb_487 : _GEN_486; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_488 = 9'h1e8 == io_ar_addr ? btb_488 : _GEN_487; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_489 = 9'h1e9 == io_ar_addr ? btb_489 : _GEN_488; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_490 = 9'h1ea == io_ar_addr ? btb_490 : _GEN_489; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_491 = 9'h1eb == io_ar_addr ? btb_491 : _GEN_490; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_492 = 9'h1ec == io_ar_addr ? btb_492 : _GEN_491; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_493 = 9'h1ed == io_ar_addr ? btb_493 : _GEN_492; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_494 = 9'h1ee == io_ar_addr ? btb_494 : _GEN_493; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_495 = 9'h1ef == io_ar_addr ? btb_495 : _GEN_494; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_496 = 9'h1f0 == io_ar_addr ? btb_496 : _GEN_495; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_497 = 9'h1f1 == io_ar_addr ? btb_497 : _GEN_496; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_498 = 9'h1f2 == io_ar_addr ? btb_498 : _GEN_497; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_499 = 9'h1f3 == io_ar_addr ? btb_499 : _GEN_498; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_500 = 9'h1f4 == io_ar_addr ? btb_500 : _GEN_499; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_501 = 9'h1f5 == io_ar_addr ? btb_501 : _GEN_500; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_502 = 9'h1f6 == io_ar_addr ? btb_502 : _GEN_501; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_503 = 9'h1f7 == io_ar_addr ? btb_503 : _GEN_502; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_504 = 9'h1f8 == io_ar_addr ? btb_504 : _GEN_503; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_505 = 9'h1f9 == io_ar_addr ? btb_505 : _GEN_504; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_506 = 9'h1fa == io_ar_addr ? btb_506 : _GEN_505; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_507 = 9'h1fb == io_ar_addr ? btb_507 : _GEN_506; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_508 = 9'h1fc == io_ar_addr ? btb_508 : _GEN_507; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_509 = 9'h1fd == io_ar_addr ? btb_509 : _GEN_508; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_510 = 9'h1fe == io_ar_addr ? btb_510 : _GEN_509; // @[ports_lookup_table.scala 82:{12,12}]
  wire [31:0] _GEN_513 = 9'h1 == io_aw_addr ? btb_1 : btb_0; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_514 = 9'h2 == io_aw_addr ? btb_2 : _GEN_513; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_515 = 9'h3 == io_aw_addr ? btb_3 : _GEN_514; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_516 = 9'h4 == io_aw_addr ? btb_4 : _GEN_515; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_517 = 9'h5 == io_aw_addr ? btb_5 : _GEN_516; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_518 = 9'h6 == io_aw_addr ? btb_6 : _GEN_517; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_519 = 9'h7 == io_aw_addr ? btb_7 : _GEN_518; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_520 = 9'h8 == io_aw_addr ? btb_8 : _GEN_519; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_521 = 9'h9 == io_aw_addr ? btb_9 : _GEN_520; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_522 = 9'ha == io_aw_addr ? btb_10 : _GEN_521; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_523 = 9'hb == io_aw_addr ? btb_11 : _GEN_522; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_524 = 9'hc == io_aw_addr ? btb_12 : _GEN_523; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_525 = 9'hd == io_aw_addr ? btb_13 : _GEN_524; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_526 = 9'he == io_aw_addr ? btb_14 : _GEN_525; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_527 = 9'hf == io_aw_addr ? btb_15 : _GEN_526; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_528 = 9'h10 == io_aw_addr ? btb_16 : _GEN_527; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_529 = 9'h11 == io_aw_addr ? btb_17 : _GEN_528; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_530 = 9'h12 == io_aw_addr ? btb_18 : _GEN_529; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_531 = 9'h13 == io_aw_addr ? btb_19 : _GEN_530; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_532 = 9'h14 == io_aw_addr ? btb_20 : _GEN_531; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_533 = 9'h15 == io_aw_addr ? btb_21 : _GEN_532; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_534 = 9'h16 == io_aw_addr ? btb_22 : _GEN_533; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_535 = 9'h17 == io_aw_addr ? btb_23 : _GEN_534; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_536 = 9'h18 == io_aw_addr ? btb_24 : _GEN_535; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_537 = 9'h19 == io_aw_addr ? btb_25 : _GEN_536; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_538 = 9'h1a == io_aw_addr ? btb_26 : _GEN_537; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_539 = 9'h1b == io_aw_addr ? btb_27 : _GEN_538; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_540 = 9'h1c == io_aw_addr ? btb_28 : _GEN_539; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_541 = 9'h1d == io_aw_addr ? btb_29 : _GEN_540; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_542 = 9'h1e == io_aw_addr ? btb_30 : _GEN_541; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_543 = 9'h1f == io_aw_addr ? btb_31 : _GEN_542; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_544 = 9'h20 == io_aw_addr ? btb_32 : _GEN_543; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_545 = 9'h21 == io_aw_addr ? btb_33 : _GEN_544; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_546 = 9'h22 == io_aw_addr ? btb_34 : _GEN_545; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_547 = 9'h23 == io_aw_addr ? btb_35 : _GEN_546; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_548 = 9'h24 == io_aw_addr ? btb_36 : _GEN_547; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_549 = 9'h25 == io_aw_addr ? btb_37 : _GEN_548; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_550 = 9'h26 == io_aw_addr ? btb_38 : _GEN_549; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_551 = 9'h27 == io_aw_addr ? btb_39 : _GEN_550; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_552 = 9'h28 == io_aw_addr ? btb_40 : _GEN_551; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_553 = 9'h29 == io_aw_addr ? btb_41 : _GEN_552; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_554 = 9'h2a == io_aw_addr ? btb_42 : _GEN_553; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_555 = 9'h2b == io_aw_addr ? btb_43 : _GEN_554; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_556 = 9'h2c == io_aw_addr ? btb_44 : _GEN_555; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_557 = 9'h2d == io_aw_addr ? btb_45 : _GEN_556; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_558 = 9'h2e == io_aw_addr ? btb_46 : _GEN_557; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_559 = 9'h2f == io_aw_addr ? btb_47 : _GEN_558; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_560 = 9'h30 == io_aw_addr ? btb_48 : _GEN_559; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_561 = 9'h31 == io_aw_addr ? btb_49 : _GEN_560; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_562 = 9'h32 == io_aw_addr ? btb_50 : _GEN_561; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_563 = 9'h33 == io_aw_addr ? btb_51 : _GEN_562; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_564 = 9'h34 == io_aw_addr ? btb_52 : _GEN_563; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_565 = 9'h35 == io_aw_addr ? btb_53 : _GEN_564; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_566 = 9'h36 == io_aw_addr ? btb_54 : _GEN_565; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_567 = 9'h37 == io_aw_addr ? btb_55 : _GEN_566; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_568 = 9'h38 == io_aw_addr ? btb_56 : _GEN_567; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_569 = 9'h39 == io_aw_addr ? btb_57 : _GEN_568; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_570 = 9'h3a == io_aw_addr ? btb_58 : _GEN_569; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_571 = 9'h3b == io_aw_addr ? btb_59 : _GEN_570; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_572 = 9'h3c == io_aw_addr ? btb_60 : _GEN_571; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_573 = 9'h3d == io_aw_addr ? btb_61 : _GEN_572; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_574 = 9'h3e == io_aw_addr ? btb_62 : _GEN_573; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_575 = 9'h3f == io_aw_addr ? btb_63 : _GEN_574; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_576 = 9'h40 == io_aw_addr ? btb_64 : _GEN_575; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_577 = 9'h41 == io_aw_addr ? btb_65 : _GEN_576; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_578 = 9'h42 == io_aw_addr ? btb_66 : _GEN_577; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_579 = 9'h43 == io_aw_addr ? btb_67 : _GEN_578; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_580 = 9'h44 == io_aw_addr ? btb_68 : _GEN_579; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_581 = 9'h45 == io_aw_addr ? btb_69 : _GEN_580; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_582 = 9'h46 == io_aw_addr ? btb_70 : _GEN_581; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_583 = 9'h47 == io_aw_addr ? btb_71 : _GEN_582; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_584 = 9'h48 == io_aw_addr ? btb_72 : _GEN_583; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_585 = 9'h49 == io_aw_addr ? btb_73 : _GEN_584; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_586 = 9'h4a == io_aw_addr ? btb_74 : _GEN_585; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_587 = 9'h4b == io_aw_addr ? btb_75 : _GEN_586; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_588 = 9'h4c == io_aw_addr ? btb_76 : _GEN_587; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_589 = 9'h4d == io_aw_addr ? btb_77 : _GEN_588; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_590 = 9'h4e == io_aw_addr ? btb_78 : _GEN_589; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_591 = 9'h4f == io_aw_addr ? btb_79 : _GEN_590; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_592 = 9'h50 == io_aw_addr ? btb_80 : _GEN_591; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_593 = 9'h51 == io_aw_addr ? btb_81 : _GEN_592; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_594 = 9'h52 == io_aw_addr ? btb_82 : _GEN_593; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_595 = 9'h53 == io_aw_addr ? btb_83 : _GEN_594; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_596 = 9'h54 == io_aw_addr ? btb_84 : _GEN_595; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_597 = 9'h55 == io_aw_addr ? btb_85 : _GEN_596; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_598 = 9'h56 == io_aw_addr ? btb_86 : _GEN_597; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_599 = 9'h57 == io_aw_addr ? btb_87 : _GEN_598; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_600 = 9'h58 == io_aw_addr ? btb_88 : _GEN_599; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_601 = 9'h59 == io_aw_addr ? btb_89 : _GEN_600; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_602 = 9'h5a == io_aw_addr ? btb_90 : _GEN_601; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_603 = 9'h5b == io_aw_addr ? btb_91 : _GEN_602; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_604 = 9'h5c == io_aw_addr ? btb_92 : _GEN_603; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_605 = 9'h5d == io_aw_addr ? btb_93 : _GEN_604; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_606 = 9'h5e == io_aw_addr ? btb_94 : _GEN_605; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_607 = 9'h5f == io_aw_addr ? btb_95 : _GEN_606; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_608 = 9'h60 == io_aw_addr ? btb_96 : _GEN_607; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_609 = 9'h61 == io_aw_addr ? btb_97 : _GEN_608; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_610 = 9'h62 == io_aw_addr ? btb_98 : _GEN_609; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_611 = 9'h63 == io_aw_addr ? btb_99 : _GEN_610; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_612 = 9'h64 == io_aw_addr ? btb_100 : _GEN_611; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_613 = 9'h65 == io_aw_addr ? btb_101 : _GEN_612; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_614 = 9'h66 == io_aw_addr ? btb_102 : _GEN_613; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_615 = 9'h67 == io_aw_addr ? btb_103 : _GEN_614; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_616 = 9'h68 == io_aw_addr ? btb_104 : _GEN_615; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_617 = 9'h69 == io_aw_addr ? btb_105 : _GEN_616; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_618 = 9'h6a == io_aw_addr ? btb_106 : _GEN_617; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_619 = 9'h6b == io_aw_addr ? btb_107 : _GEN_618; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_620 = 9'h6c == io_aw_addr ? btb_108 : _GEN_619; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_621 = 9'h6d == io_aw_addr ? btb_109 : _GEN_620; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_622 = 9'h6e == io_aw_addr ? btb_110 : _GEN_621; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_623 = 9'h6f == io_aw_addr ? btb_111 : _GEN_622; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_624 = 9'h70 == io_aw_addr ? btb_112 : _GEN_623; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_625 = 9'h71 == io_aw_addr ? btb_113 : _GEN_624; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_626 = 9'h72 == io_aw_addr ? btb_114 : _GEN_625; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_627 = 9'h73 == io_aw_addr ? btb_115 : _GEN_626; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_628 = 9'h74 == io_aw_addr ? btb_116 : _GEN_627; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_629 = 9'h75 == io_aw_addr ? btb_117 : _GEN_628; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_630 = 9'h76 == io_aw_addr ? btb_118 : _GEN_629; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_631 = 9'h77 == io_aw_addr ? btb_119 : _GEN_630; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_632 = 9'h78 == io_aw_addr ? btb_120 : _GEN_631; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_633 = 9'h79 == io_aw_addr ? btb_121 : _GEN_632; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_634 = 9'h7a == io_aw_addr ? btb_122 : _GEN_633; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_635 = 9'h7b == io_aw_addr ? btb_123 : _GEN_634; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_636 = 9'h7c == io_aw_addr ? btb_124 : _GEN_635; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_637 = 9'h7d == io_aw_addr ? btb_125 : _GEN_636; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_638 = 9'h7e == io_aw_addr ? btb_126 : _GEN_637; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_639 = 9'h7f == io_aw_addr ? btb_127 : _GEN_638; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_640 = 9'h80 == io_aw_addr ? btb_128 : _GEN_639; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_641 = 9'h81 == io_aw_addr ? btb_129 : _GEN_640; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_642 = 9'h82 == io_aw_addr ? btb_130 : _GEN_641; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_643 = 9'h83 == io_aw_addr ? btb_131 : _GEN_642; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_644 = 9'h84 == io_aw_addr ? btb_132 : _GEN_643; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_645 = 9'h85 == io_aw_addr ? btb_133 : _GEN_644; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_646 = 9'h86 == io_aw_addr ? btb_134 : _GEN_645; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_647 = 9'h87 == io_aw_addr ? btb_135 : _GEN_646; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_648 = 9'h88 == io_aw_addr ? btb_136 : _GEN_647; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_649 = 9'h89 == io_aw_addr ? btb_137 : _GEN_648; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_650 = 9'h8a == io_aw_addr ? btb_138 : _GEN_649; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_651 = 9'h8b == io_aw_addr ? btb_139 : _GEN_650; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_652 = 9'h8c == io_aw_addr ? btb_140 : _GEN_651; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_653 = 9'h8d == io_aw_addr ? btb_141 : _GEN_652; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_654 = 9'h8e == io_aw_addr ? btb_142 : _GEN_653; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_655 = 9'h8f == io_aw_addr ? btb_143 : _GEN_654; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_656 = 9'h90 == io_aw_addr ? btb_144 : _GEN_655; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_657 = 9'h91 == io_aw_addr ? btb_145 : _GEN_656; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_658 = 9'h92 == io_aw_addr ? btb_146 : _GEN_657; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_659 = 9'h93 == io_aw_addr ? btb_147 : _GEN_658; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_660 = 9'h94 == io_aw_addr ? btb_148 : _GEN_659; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_661 = 9'h95 == io_aw_addr ? btb_149 : _GEN_660; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_662 = 9'h96 == io_aw_addr ? btb_150 : _GEN_661; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_663 = 9'h97 == io_aw_addr ? btb_151 : _GEN_662; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_664 = 9'h98 == io_aw_addr ? btb_152 : _GEN_663; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_665 = 9'h99 == io_aw_addr ? btb_153 : _GEN_664; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_666 = 9'h9a == io_aw_addr ? btb_154 : _GEN_665; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_667 = 9'h9b == io_aw_addr ? btb_155 : _GEN_666; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_668 = 9'h9c == io_aw_addr ? btb_156 : _GEN_667; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_669 = 9'h9d == io_aw_addr ? btb_157 : _GEN_668; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_670 = 9'h9e == io_aw_addr ? btb_158 : _GEN_669; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_671 = 9'h9f == io_aw_addr ? btb_159 : _GEN_670; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_672 = 9'ha0 == io_aw_addr ? btb_160 : _GEN_671; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_673 = 9'ha1 == io_aw_addr ? btb_161 : _GEN_672; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_674 = 9'ha2 == io_aw_addr ? btb_162 : _GEN_673; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_675 = 9'ha3 == io_aw_addr ? btb_163 : _GEN_674; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_676 = 9'ha4 == io_aw_addr ? btb_164 : _GEN_675; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_677 = 9'ha5 == io_aw_addr ? btb_165 : _GEN_676; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_678 = 9'ha6 == io_aw_addr ? btb_166 : _GEN_677; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_679 = 9'ha7 == io_aw_addr ? btb_167 : _GEN_678; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_680 = 9'ha8 == io_aw_addr ? btb_168 : _GEN_679; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_681 = 9'ha9 == io_aw_addr ? btb_169 : _GEN_680; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_682 = 9'haa == io_aw_addr ? btb_170 : _GEN_681; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_683 = 9'hab == io_aw_addr ? btb_171 : _GEN_682; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_684 = 9'hac == io_aw_addr ? btb_172 : _GEN_683; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_685 = 9'had == io_aw_addr ? btb_173 : _GEN_684; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_686 = 9'hae == io_aw_addr ? btb_174 : _GEN_685; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_687 = 9'haf == io_aw_addr ? btb_175 : _GEN_686; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_688 = 9'hb0 == io_aw_addr ? btb_176 : _GEN_687; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_689 = 9'hb1 == io_aw_addr ? btb_177 : _GEN_688; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_690 = 9'hb2 == io_aw_addr ? btb_178 : _GEN_689; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_691 = 9'hb3 == io_aw_addr ? btb_179 : _GEN_690; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_692 = 9'hb4 == io_aw_addr ? btb_180 : _GEN_691; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_693 = 9'hb5 == io_aw_addr ? btb_181 : _GEN_692; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_694 = 9'hb6 == io_aw_addr ? btb_182 : _GEN_693; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_695 = 9'hb7 == io_aw_addr ? btb_183 : _GEN_694; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_696 = 9'hb8 == io_aw_addr ? btb_184 : _GEN_695; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_697 = 9'hb9 == io_aw_addr ? btb_185 : _GEN_696; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_698 = 9'hba == io_aw_addr ? btb_186 : _GEN_697; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_699 = 9'hbb == io_aw_addr ? btb_187 : _GEN_698; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_700 = 9'hbc == io_aw_addr ? btb_188 : _GEN_699; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_701 = 9'hbd == io_aw_addr ? btb_189 : _GEN_700; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_702 = 9'hbe == io_aw_addr ? btb_190 : _GEN_701; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_703 = 9'hbf == io_aw_addr ? btb_191 : _GEN_702; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_704 = 9'hc0 == io_aw_addr ? btb_192 : _GEN_703; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_705 = 9'hc1 == io_aw_addr ? btb_193 : _GEN_704; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_706 = 9'hc2 == io_aw_addr ? btb_194 : _GEN_705; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_707 = 9'hc3 == io_aw_addr ? btb_195 : _GEN_706; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_708 = 9'hc4 == io_aw_addr ? btb_196 : _GEN_707; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_709 = 9'hc5 == io_aw_addr ? btb_197 : _GEN_708; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_710 = 9'hc6 == io_aw_addr ? btb_198 : _GEN_709; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_711 = 9'hc7 == io_aw_addr ? btb_199 : _GEN_710; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_712 = 9'hc8 == io_aw_addr ? btb_200 : _GEN_711; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_713 = 9'hc9 == io_aw_addr ? btb_201 : _GEN_712; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_714 = 9'hca == io_aw_addr ? btb_202 : _GEN_713; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_715 = 9'hcb == io_aw_addr ? btb_203 : _GEN_714; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_716 = 9'hcc == io_aw_addr ? btb_204 : _GEN_715; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_717 = 9'hcd == io_aw_addr ? btb_205 : _GEN_716; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_718 = 9'hce == io_aw_addr ? btb_206 : _GEN_717; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_719 = 9'hcf == io_aw_addr ? btb_207 : _GEN_718; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_720 = 9'hd0 == io_aw_addr ? btb_208 : _GEN_719; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_721 = 9'hd1 == io_aw_addr ? btb_209 : _GEN_720; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_722 = 9'hd2 == io_aw_addr ? btb_210 : _GEN_721; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_723 = 9'hd3 == io_aw_addr ? btb_211 : _GEN_722; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_724 = 9'hd4 == io_aw_addr ? btb_212 : _GEN_723; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_725 = 9'hd5 == io_aw_addr ? btb_213 : _GEN_724; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_726 = 9'hd6 == io_aw_addr ? btb_214 : _GEN_725; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_727 = 9'hd7 == io_aw_addr ? btb_215 : _GEN_726; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_728 = 9'hd8 == io_aw_addr ? btb_216 : _GEN_727; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_729 = 9'hd9 == io_aw_addr ? btb_217 : _GEN_728; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_730 = 9'hda == io_aw_addr ? btb_218 : _GEN_729; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_731 = 9'hdb == io_aw_addr ? btb_219 : _GEN_730; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_732 = 9'hdc == io_aw_addr ? btb_220 : _GEN_731; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_733 = 9'hdd == io_aw_addr ? btb_221 : _GEN_732; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_734 = 9'hde == io_aw_addr ? btb_222 : _GEN_733; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_735 = 9'hdf == io_aw_addr ? btb_223 : _GEN_734; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_736 = 9'he0 == io_aw_addr ? btb_224 : _GEN_735; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_737 = 9'he1 == io_aw_addr ? btb_225 : _GEN_736; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_738 = 9'he2 == io_aw_addr ? btb_226 : _GEN_737; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_739 = 9'he3 == io_aw_addr ? btb_227 : _GEN_738; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_740 = 9'he4 == io_aw_addr ? btb_228 : _GEN_739; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_741 = 9'he5 == io_aw_addr ? btb_229 : _GEN_740; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_742 = 9'he6 == io_aw_addr ? btb_230 : _GEN_741; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_743 = 9'he7 == io_aw_addr ? btb_231 : _GEN_742; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_744 = 9'he8 == io_aw_addr ? btb_232 : _GEN_743; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_745 = 9'he9 == io_aw_addr ? btb_233 : _GEN_744; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_746 = 9'hea == io_aw_addr ? btb_234 : _GEN_745; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_747 = 9'heb == io_aw_addr ? btb_235 : _GEN_746; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_748 = 9'hec == io_aw_addr ? btb_236 : _GEN_747; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_749 = 9'hed == io_aw_addr ? btb_237 : _GEN_748; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_750 = 9'hee == io_aw_addr ? btb_238 : _GEN_749; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_751 = 9'hef == io_aw_addr ? btb_239 : _GEN_750; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_752 = 9'hf0 == io_aw_addr ? btb_240 : _GEN_751; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_753 = 9'hf1 == io_aw_addr ? btb_241 : _GEN_752; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_754 = 9'hf2 == io_aw_addr ? btb_242 : _GEN_753; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_755 = 9'hf3 == io_aw_addr ? btb_243 : _GEN_754; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_756 = 9'hf4 == io_aw_addr ? btb_244 : _GEN_755; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_757 = 9'hf5 == io_aw_addr ? btb_245 : _GEN_756; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_758 = 9'hf6 == io_aw_addr ? btb_246 : _GEN_757; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_759 = 9'hf7 == io_aw_addr ? btb_247 : _GEN_758; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_760 = 9'hf8 == io_aw_addr ? btb_248 : _GEN_759; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_761 = 9'hf9 == io_aw_addr ? btb_249 : _GEN_760; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_762 = 9'hfa == io_aw_addr ? btb_250 : _GEN_761; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_763 = 9'hfb == io_aw_addr ? btb_251 : _GEN_762; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_764 = 9'hfc == io_aw_addr ? btb_252 : _GEN_763; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_765 = 9'hfd == io_aw_addr ? btb_253 : _GEN_764; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_766 = 9'hfe == io_aw_addr ? btb_254 : _GEN_765; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_767 = 9'hff == io_aw_addr ? btb_255 : _GEN_766; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_768 = 9'h100 == io_aw_addr ? btb_256 : _GEN_767; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_769 = 9'h101 == io_aw_addr ? btb_257 : _GEN_768; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_770 = 9'h102 == io_aw_addr ? btb_258 : _GEN_769; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_771 = 9'h103 == io_aw_addr ? btb_259 : _GEN_770; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_772 = 9'h104 == io_aw_addr ? btb_260 : _GEN_771; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_773 = 9'h105 == io_aw_addr ? btb_261 : _GEN_772; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_774 = 9'h106 == io_aw_addr ? btb_262 : _GEN_773; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_775 = 9'h107 == io_aw_addr ? btb_263 : _GEN_774; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_776 = 9'h108 == io_aw_addr ? btb_264 : _GEN_775; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_777 = 9'h109 == io_aw_addr ? btb_265 : _GEN_776; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_778 = 9'h10a == io_aw_addr ? btb_266 : _GEN_777; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_779 = 9'h10b == io_aw_addr ? btb_267 : _GEN_778; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_780 = 9'h10c == io_aw_addr ? btb_268 : _GEN_779; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_781 = 9'h10d == io_aw_addr ? btb_269 : _GEN_780; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_782 = 9'h10e == io_aw_addr ? btb_270 : _GEN_781; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_783 = 9'h10f == io_aw_addr ? btb_271 : _GEN_782; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_784 = 9'h110 == io_aw_addr ? btb_272 : _GEN_783; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_785 = 9'h111 == io_aw_addr ? btb_273 : _GEN_784; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_786 = 9'h112 == io_aw_addr ? btb_274 : _GEN_785; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_787 = 9'h113 == io_aw_addr ? btb_275 : _GEN_786; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_788 = 9'h114 == io_aw_addr ? btb_276 : _GEN_787; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_789 = 9'h115 == io_aw_addr ? btb_277 : _GEN_788; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_790 = 9'h116 == io_aw_addr ? btb_278 : _GEN_789; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_791 = 9'h117 == io_aw_addr ? btb_279 : _GEN_790; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_792 = 9'h118 == io_aw_addr ? btb_280 : _GEN_791; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_793 = 9'h119 == io_aw_addr ? btb_281 : _GEN_792; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_794 = 9'h11a == io_aw_addr ? btb_282 : _GEN_793; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_795 = 9'h11b == io_aw_addr ? btb_283 : _GEN_794; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_796 = 9'h11c == io_aw_addr ? btb_284 : _GEN_795; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_797 = 9'h11d == io_aw_addr ? btb_285 : _GEN_796; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_798 = 9'h11e == io_aw_addr ? btb_286 : _GEN_797; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_799 = 9'h11f == io_aw_addr ? btb_287 : _GEN_798; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_800 = 9'h120 == io_aw_addr ? btb_288 : _GEN_799; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_801 = 9'h121 == io_aw_addr ? btb_289 : _GEN_800; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_802 = 9'h122 == io_aw_addr ? btb_290 : _GEN_801; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_803 = 9'h123 == io_aw_addr ? btb_291 : _GEN_802; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_804 = 9'h124 == io_aw_addr ? btb_292 : _GEN_803; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_805 = 9'h125 == io_aw_addr ? btb_293 : _GEN_804; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_806 = 9'h126 == io_aw_addr ? btb_294 : _GEN_805; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_807 = 9'h127 == io_aw_addr ? btb_295 : _GEN_806; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_808 = 9'h128 == io_aw_addr ? btb_296 : _GEN_807; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_809 = 9'h129 == io_aw_addr ? btb_297 : _GEN_808; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_810 = 9'h12a == io_aw_addr ? btb_298 : _GEN_809; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_811 = 9'h12b == io_aw_addr ? btb_299 : _GEN_810; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_812 = 9'h12c == io_aw_addr ? btb_300 : _GEN_811; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_813 = 9'h12d == io_aw_addr ? btb_301 : _GEN_812; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_814 = 9'h12e == io_aw_addr ? btb_302 : _GEN_813; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_815 = 9'h12f == io_aw_addr ? btb_303 : _GEN_814; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_816 = 9'h130 == io_aw_addr ? btb_304 : _GEN_815; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_817 = 9'h131 == io_aw_addr ? btb_305 : _GEN_816; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_818 = 9'h132 == io_aw_addr ? btb_306 : _GEN_817; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_819 = 9'h133 == io_aw_addr ? btb_307 : _GEN_818; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_820 = 9'h134 == io_aw_addr ? btb_308 : _GEN_819; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_821 = 9'h135 == io_aw_addr ? btb_309 : _GEN_820; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_822 = 9'h136 == io_aw_addr ? btb_310 : _GEN_821; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_823 = 9'h137 == io_aw_addr ? btb_311 : _GEN_822; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_824 = 9'h138 == io_aw_addr ? btb_312 : _GEN_823; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_825 = 9'h139 == io_aw_addr ? btb_313 : _GEN_824; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_826 = 9'h13a == io_aw_addr ? btb_314 : _GEN_825; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_827 = 9'h13b == io_aw_addr ? btb_315 : _GEN_826; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_828 = 9'h13c == io_aw_addr ? btb_316 : _GEN_827; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_829 = 9'h13d == io_aw_addr ? btb_317 : _GEN_828; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_830 = 9'h13e == io_aw_addr ? btb_318 : _GEN_829; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_831 = 9'h13f == io_aw_addr ? btb_319 : _GEN_830; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_832 = 9'h140 == io_aw_addr ? btb_320 : _GEN_831; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_833 = 9'h141 == io_aw_addr ? btb_321 : _GEN_832; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_834 = 9'h142 == io_aw_addr ? btb_322 : _GEN_833; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_835 = 9'h143 == io_aw_addr ? btb_323 : _GEN_834; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_836 = 9'h144 == io_aw_addr ? btb_324 : _GEN_835; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_837 = 9'h145 == io_aw_addr ? btb_325 : _GEN_836; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_838 = 9'h146 == io_aw_addr ? btb_326 : _GEN_837; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_839 = 9'h147 == io_aw_addr ? btb_327 : _GEN_838; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_840 = 9'h148 == io_aw_addr ? btb_328 : _GEN_839; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_841 = 9'h149 == io_aw_addr ? btb_329 : _GEN_840; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_842 = 9'h14a == io_aw_addr ? btb_330 : _GEN_841; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_843 = 9'h14b == io_aw_addr ? btb_331 : _GEN_842; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_844 = 9'h14c == io_aw_addr ? btb_332 : _GEN_843; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_845 = 9'h14d == io_aw_addr ? btb_333 : _GEN_844; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_846 = 9'h14e == io_aw_addr ? btb_334 : _GEN_845; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_847 = 9'h14f == io_aw_addr ? btb_335 : _GEN_846; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_848 = 9'h150 == io_aw_addr ? btb_336 : _GEN_847; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_849 = 9'h151 == io_aw_addr ? btb_337 : _GEN_848; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_850 = 9'h152 == io_aw_addr ? btb_338 : _GEN_849; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_851 = 9'h153 == io_aw_addr ? btb_339 : _GEN_850; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_852 = 9'h154 == io_aw_addr ? btb_340 : _GEN_851; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_853 = 9'h155 == io_aw_addr ? btb_341 : _GEN_852; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_854 = 9'h156 == io_aw_addr ? btb_342 : _GEN_853; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_855 = 9'h157 == io_aw_addr ? btb_343 : _GEN_854; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_856 = 9'h158 == io_aw_addr ? btb_344 : _GEN_855; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_857 = 9'h159 == io_aw_addr ? btb_345 : _GEN_856; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_858 = 9'h15a == io_aw_addr ? btb_346 : _GEN_857; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_859 = 9'h15b == io_aw_addr ? btb_347 : _GEN_858; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_860 = 9'h15c == io_aw_addr ? btb_348 : _GEN_859; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_861 = 9'h15d == io_aw_addr ? btb_349 : _GEN_860; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_862 = 9'h15e == io_aw_addr ? btb_350 : _GEN_861; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_863 = 9'h15f == io_aw_addr ? btb_351 : _GEN_862; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_864 = 9'h160 == io_aw_addr ? btb_352 : _GEN_863; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_865 = 9'h161 == io_aw_addr ? btb_353 : _GEN_864; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_866 = 9'h162 == io_aw_addr ? btb_354 : _GEN_865; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_867 = 9'h163 == io_aw_addr ? btb_355 : _GEN_866; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_868 = 9'h164 == io_aw_addr ? btb_356 : _GEN_867; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_869 = 9'h165 == io_aw_addr ? btb_357 : _GEN_868; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_870 = 9'h166 == io_aw_addr ? btb_358 : _GEN_869; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_871 = 9'h167 == io_aw_addr ? btb_359 : _GEN_870; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_872 = 9'h168 == io_aw_addr ? btb_360 : _GEN_871; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_873 = 9'h169 == io_aw_addr ? btb_361 : _GEN_872; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_874 = 9'h16a == io_aw_addr ? btb_362 : _GEN_873; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_875 = 9'h16b == io_aw_addr ? btb_363 : _GEN_874; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_876 = 9'h16c == io_aw_addr ? btb_364 : _GEN_875; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_877 = 9'h16d == io_aw_addr ? btb_365 : _GEN_876; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_878 = 9'h16e == io_aw_addr ? btb_366 : _GEN_877; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_879 = 9'h16f == io_aw_addr ? btb_367 : _GEN_878; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_880 = 9'h170 == io_aw_addr ? btb_368 : _GEN_879; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_881 = 9'h171 == io_aw_addr ? btb_369 : _GEN_880; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_882 = 9'h172 == io_aw_addr ? btb_370 : _GEN_881; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_883 = 9'h173 == io_aw_addr ? btb_371 : _GEN_882; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_884 = 9'h174 == io_aw_addr ? btb_372 : _GEN_883; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_885 = 9'h175 == io_aw_addr ? btb_373 : _GEN_884; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_886 = 9'h176 == io_aw_addr ? btb_374 : _GEN_885; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_887 = 9'h177 == io_aw_addr ? btb_375 : _GEN_886; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_888 = 9'h178 == io_aw_addr ? btb_376 : _GEN_887; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_889 = 9'h179 == io_aw_addr ? btb_377 : _GEN_888; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_890 = 9'h17a == io_aw_addr ? btb_378 : _GEN_889; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_891 = 9'h17b == io_aw_addr ? btb_379 : _GEN_890; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_892 = 9'h17c == io_aw_addr ? btb_380 : _GEN_891; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_893 = 9'h17d == io_aw_addr ? btb_381 : _GEN_892; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_894 = 9'h17e == io_aw_addr ? btb_382 : _GEN_893; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_895 = 9'h17f == io_aw_addr ? btb_383 : _GEN_894; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_896 = 9'h180 == io_aw_addr ? btb_384 : _GEN_895; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_897 = 9'h181 == io_aw_addr ? btb_385 : _GEN_896; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_898 = 9'h182 == io_aw_addr ? btb_386 : _GEN_897; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_899 = 9'h183 == io_aw_addr ? btb_387 : _GEN_898; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_900 = 9'h184 == io_aw_addr ? btb_388 : _GEN_899; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_901 = 9'h185 == io_aw_addr ? btb_389 : _GEN_900; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_902 = 9'h186 == io_aw_addr ? btb_390 : _GEN_901; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_903 = 9'h187 == io_aw_addr ? btb_391 : _GEN_902; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_904 = 9'h188 == io_aw_addr ? btb_392 : _GEN_903; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_905 = 9'h189 == io_aw_addr ? btb_393 : _GEN_904; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_906 = 9'h18a == io_aw_addr ? btb_394 : _GEN_905; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_907 = 9'h18b == io_aw_addr ? btb_395 : _GEN_906; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_908 = 9'h18c == io_aw_addr ? btb_396 : _GEN_907; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_909 = 9'h18d == io_aw_addr ? btb_397 : _GEN_908; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_910 = 9'h18e == io_aw_addr ? btb_398 : _GEN_909; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_911 = 9'h18f == io_aw_addr ? btb_399 : _GEN_910; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_912 = 9'h190 == io_aw_addr ? btb_400 : _GEN_911; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_913 = 9'h191 == io_aw_addr ? btb_401 : _GEN_912; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_914 = 9'h192 == io_aw_addr ? btb_402 : _GEN_913; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_915 = 9'h193 == io_aw_addr ? btb_403 : _GEN_914; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_916 = 9'h194 == io_aw_addr ? btb_404 : _GEN_915; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_917 = 9'h195 == io_aw_addr ? btb_405 : _GEN_916; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_918 = 9'h196 == io_aw_addr ? btb_406 : _GEN_917; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_919 = 9'h197 == io_aw_addr ? btb_407 : _GEN_918; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_920 = 9'h198 == io_aw_addr ? btb_408 : _GEN_919; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_921 = 9'h199 == io_aw_addr ? btb_409 : _GEN_920; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_922 = 9'h19a == io_aw_addr ? btb_410 : _GEN_921; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_923 = 9'h19b == io_aw_addr ? btb_411 : _GEN_922; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_924 = 9'h19c == io_aw_addr ? btb_412 : _GEN_923; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_925 = 9'h19d == io_aw_addr ? btb_413 : _GEN_924; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_926 = 9'h19e == io_aw_addr ? btb_414 : _GEN_925; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_927 = 9'h19f == io_aw_addr ? btb_415 : _GEN_926; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_928 = 9'h1a0 == io_aw_addr ? btb_416 : _GEN_927; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_929 = 9'h1a1 == io_aw_addr ? btb_417 : _GEN_928; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_930 = 9'h1a2 == io_aw_addr ? btb_418 : _GEN_929; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_931 = 9'h1a3 == io_aw_addr ? btb_419 : _GEN_930; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_932 = 9'h1a4 == io_aw_addr ? btb_420 : _GEN_931; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_933 = 9'h1a5 == io_aw_addr ? btb_421 : _GEN_932; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_934 = 9'h1a6 == io_aw_addr ? btb_422 : _GEN_933; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_935 = 9'h1a7 == io_aw_addr ? btb_423 : _GEN_934; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_936 = 9'h1a8 == io_aw_addr ? btb_424 : _GEN_935; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_937 = 9'h1a9 == io_aw_addr ? btb_425 : _GEN_936; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_938 = 9'h1aa == io_aw_addr ? btb_426 : _GEN_937; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_939 = 9'h1ab == io_aw_addr ? btb_427 : _GEN_938; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_940 = 9'h1ac == io_aw_addr ? btb_428 : _GEN_939; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_941 = 9'h1ad == io_aw_addr ? btb_429 : _GEN_940; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_942 = 9'h1ae == io_aw_addr ? btb_430 : _GEN_941; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_943 = 9'h1af == io_aw_addr ? btb_431 : _GEN_942; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_944 = 9'h1b0 == io_aw_addr ? btb_432 : _GEN_943; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_945 = 9'h1b1 == io_aw_addr ? btb_433 : _GEN_944; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_946 = 9'h1b2 == io_aw_addr ? btb_434 : _GEN_945; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_947 = 9'h1b3 == io_aw_addr ? btb_435 : _GEN_946; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_948 = 9'h1b4 == io_aw_addr ? btb_436 : _GEN_947; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_949 = 9'h1b5 == io_aw_addr ? btb_437 : _GEN_948; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_950 = 9'h1b6 == io_aw_addr ? btb_438 : _GEN_949; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_951 = 9'h1b7 == io_aw_addr ? btb_439 : _GEN_950; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_952 = 9'h1b8 == io_aw_addr ? btb_440 : _GEN_951; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_953 = 9'h1b9 == io_aw_addr ? btb_441 : _GEN_952; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_954 = 9'h1ba == io_aw_addr ? btb_442 : _GEN_953; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_955 = 9'h1bb == io_aw_addr ? btb_443 : _GEN_954; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_956 = 9'h1bc == io_aw_addr ? btb_444 : _GEN_955; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_957 = 9'h1bd == io_aw_addr ? btb_445 : _GEN_956; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_958 = 9'h1be == io_aw_addr ? btb_446 : _GEN_957; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_959 = 9'h1bf == io_aw_addr ? btb_447 : _GEN_958; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_960 = 9'h1c0 == io_aw_addr ? btb_448 : _GEN_959; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_961 = 9'h1c1 == io_aw_addr ? btb_449 : _GEN_960; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_962 = 9'h1c2 == io_aw_addr ? btb_450 : _GEN_961; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_963 = 9'h1c3 == io_aw_addr ? btb_451 : _GEN_962; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_964 = 9'h1c4 == io_aw_addr ? btb_452 : _GEN_963; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_965 = 9'h1c5 == io_aw_addr ? btb_453 : _GEN_964; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_966 = 9'h1c6 == io_aw_addr ? btb_454 : _GEN_965; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_967 = 9'h1c7 == io_aw_addr ? btb_455 : _GEN_966; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_968 = 9'h1c8 == io_aw_addr ? btb_456 : _GEN_967; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_969 = 9'h1c9 == io_aw_addr ? btb_457 : _GEN_968; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_970 = 9'h1ca == io_aw_addr ? btb_458 : _GEN_969; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_971 = 9'h1cb == io_aw_addr ? btb_459 : _GEN_970; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_972 = 9'h1cc == io_aw_addr ? btb_460 : _GEN_971; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_973 = 9'h1cd == io_aw_addr ? btb_461 : _GEN_972; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_974 = 9'h1ce == io_aw_addr ? btb_462 : _GEN_973; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_975 = 9'h1cf == io_aw_addr ? btb_463 : _GEN_974; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_976 = 9'h1d0 == io_aw_addr ? btb_464 : _GEN_975; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_977 = 9'h1d1 == io_aw_addr ? btb_465 : _GEN_976; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_978 = 9'h1d2 == io_aw_addr ? btb_466 : _GEN_977; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_979 = 9'h1d3 == io_aw_addr ? btb_467 : _GEN_978; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_980 = 9'h1d4 == io_aw_addr ? btb_468 : _GEN_979; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_981 = 9'h1d5 == io_aw_addr ? btb_469 : _GEN_980; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_982 = 9'h1d6 == io_aw_addr ? btb_470 : _GEN_981; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_983 = 9'h1d7 == io_aw_addr ? btb_471 : _GEN_982; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_984 = 9'h1d8 == io_aw_addr ? btb_472 : _GEN_983; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_985 = 9'h1d9 == io_aw_addr ? btb_473 : _GEN_984; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_986 = 9'h1da == io_aw_addr ? btb_474 : _GEN_985; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_987 = 9'h1db == io_aw_addr ? btb_475 : _GEN_986; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_988 = 9'h1dc == io_aw_addr ? btb_476 : _GEN_987; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_989 = 9'h1dd == io_aw_addr ? btb_477 : _GEN_988; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_990 = 9'h1de == io_aw_addr ? btb_478 : _GEN_989; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_991 = 9'h1df == io_aw_addr ? btb_479 : _GEN_990; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_992 = 9'h1e0 == io_aw_addr ? btb_480 : _GEN_991; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_993 = 9'h1e1 == io_aw_addr ? btb_481 : _GEN_992; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_994 = 9'h1e2 == io_aw_addr ? btb_482 : _GEN_993; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_995 = 9'h1e3 == io_aw_addr ? btb_483 : _GEN_994; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_996 = 9'h1e4 == io_aw_addr ? btb_484 : _GEN_995; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_997 = 9'h1e5 == io_aw_addr ? btb_485 : _GEN_996; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_998 = 9'h1e6 == io_aw_addr ? btb_486 : _GEN_997; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_999 = 9'h1e7 == io_aw_addr ? btb_487 : _GEN_998; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1000 = 9'h1e8 == io_aw_addr ? btb_488 : _GEN_999; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1001 = 9'h1e9 == io_aw_addr ? btb_489 : _GEN_1000; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1002 = 9'h1ea == io_aw_addr ? btb_490 : _GEN_1001; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1003 = 9'h1eb == io_aw_addr ? btb_491 : _GEN_1002; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1004 = 9'h1ec == io_aw_addr ? btb_492 : _GEN_1003; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1005 = 9'h1ed == io_aw_addr ? btb_493 : _GEN_1004; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1006 = 9'h1ee == io_aw_addr ? btb_494 : _GEN_1005; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1007 = 9'h1ef == io_aw_addr ? btb_495 : _GEN_1006; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1008 = 9'h1f0 == io_aw_addr ? btb_496 : _GEN_1007; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1009 = 9'h1f1 == io_aw_addr ? btb_497 : _GEN_1008; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1010 = 9'h1f2 == io_aw_addr ? btb_498 : _GEN_1009; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1011 = 9'h1f3 == io_aw_addr ? btb_499 : _GEN_1010; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1012 = 9'h1f4 == io_aw_addr ? btb_500 : _GEN_1011; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1013 = 9'h1f5 == io_aw_addr ? btb_501 : _GEN_1012; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1014 = 9'h1f6 == io_aw_addr ? btb_502 : _GEN_1013; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1015 = 9'h1f7 == io_aw_addr ? btb_503 : _GEN_1014; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1016 = 9'h1f8 == io_aw_addr ? btb_504 : _GEN_1015; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1017 = 9'h1f9 == io_aw_addr ? btb_505 : _GEN_1016; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1018 = 9'h1fa == io_aw_addr ? btb_506 : _GEN_1017; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1019 = 9'h1fb == io_aw_addr ? btb_507 : _GEN_1018; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1020 = 9'h1fc == io_aw_addr ? btb_508 : _GEN_1019; // @[ports_lookup_table.scala 83:{27,27}]
  wire [31:0] _GEN_1021 = 9'h1fd == io_aw_addr ? btb_509 : _GEN_1020; // @[ports_lookup_table.scala 83:{27,27}]
  assign io_out = 9'h1ff == io_ar_addr ? btb_511 : _GEN_510; // @[ports_lookup_table.scala 82:{12,12}]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_0 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_0 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_0 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_0 <= btb_510;
      end else begin
        btb_0 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_1 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_1 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_1 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_1 <= btb_510;
      end else begin
        btb_1 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_2 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_2 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_2 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_2 <= btb_510;
      end else begin
        btb_2 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_3 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_3 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_3 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_3 <= btb_510;
      end else begin
        btb_3 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_4 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_4 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_4 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_4 <= btb_510;
      end else begin
        btb_4 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_5 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_5 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_5 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_5 <= btb_510;
      end else begin
        btb_5 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_6 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_6 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_6 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_6 <= btb_510;
      end else begin
        btb_6 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_7 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_7 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_7 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_7 <= btb_510;
      end else begin
        btb_7 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_8 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_8 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_8 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_8 <= btb_510;
      end else begin
        btb_8 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_9 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_9 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_9 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_9 <= btb_510;
      end else begin
        btb_9 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_10 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_10 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_10 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_10 <= btb_510;
      end else begin
        btb_10 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_11 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_11 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_11 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_11 <= btb_510;
      end else begin
        btb_11 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_12 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_12 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_12 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_12 <= btb_510;
      end else begin
        btb_12 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_13 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_13 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_13 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_13 <= btb_510;
      end else begin
        btb_13 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_14 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_14 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_14 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_14 <= btb_510;
      end else begin
        btb_14 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_15 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_15 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_15 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_15 <= btb_510;
      end else begin
        btb_15 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_16 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h10 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_16 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_16 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_16 <= btb_510;
      end else begin
        btb_16 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_17 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h11 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_17 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_17 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_17 <= btb_510;
      end else begin
        btb_17 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_18 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h12 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_18 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_18 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_18 <= btb_510;
      end else begin
        btb_18 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_19 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h13 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_19 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_19 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_19 <= btb_510;
      end else begin
        btb_19 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_20 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h14 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_20 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_20 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_20 <= btb_510;
      end else begin
        btb_20 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_21 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h15 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_21 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_21 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_21 <= btb_510;
      end else begin
        btb_21 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_22 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h16 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_22 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_22 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_22 <= btb_510;
      end else begin
        btb_22 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_23 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h17 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_23 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_23 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_23 <= btb_510;
      end else begin
        btb_23 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_24 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h18 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_24 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_24 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_24 <= btb_510;
      end else begin
        btb_24 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_25 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h19 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_25 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_25 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_25 <= btb_510;
      end else begin
        btb_25 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_26 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_26 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_26 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_26 <= btb_510;
      end else begin
        btb_26 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_27 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_27 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_27 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_27 <= btb_510;
      end else begin
        btb_27 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_28 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_28 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_28 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_28 <= btb_510;
      end else begin
        btb_28 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_29 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_29 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_29 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_29 <= btb_510;
      end else begin
        btb_29 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_30 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_30 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_30 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_30 <= btb_510;
      end else begin
        btb_30 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_31 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_31 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_31 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_31 <= btb_510;
      end else begin
        btb_31 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_32 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h20 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_32 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_32 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_32 <= btb_510;
      end else begin
        btb_32 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_33 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h21 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_33 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_33 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_33 <= btb_510;
      end else begin
        btb_33 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_34 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h22 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_34 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_34 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_34 <= btb_510;
      end else begin
        btb_34 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_35 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h23 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_35 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_35 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_35 <= btb_510;
      end else begin
        btb_35 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_36 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h24 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_36 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_36 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_36 <= btb_510;
      end else begin
        btb_36 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_37 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h25 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_37 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_37 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_37 <= btb_510;
      end else begin
        btb_37 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_38 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h26 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_38 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_38 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_38 <= btb_510;
      end else begin
        btb_38 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_39 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h27 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_39 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_39 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_39 <= btb_510;
      end else begin
        btb_39 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_40 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h28 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_40 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_40 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_40 <= btb_510;
      end else begin
        btb_40 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_41 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h29 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_41 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_41 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_41 <= btb_510;
      end else begin
        btb_41 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_42 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h2a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_42 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_42 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_42 <= btb_510;
      end else begin
        btb_42 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_43 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h2b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_43 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_43 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_43 <= btb_510;
      end else begin
        btb_43 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_44 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h2c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_44 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_44 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_44 <= btb_510;
      end else begin
        btb_44 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_45 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h2d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_45 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_45 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_45 <= btb_510;
      end else begin
        btb_45 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_46 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h2e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_46 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_46 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_46 <= btb_510;
      end else begin
        btb_46 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_47 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h2f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_47 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_47 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_47 <= btb_510;
      end else begin
        btb_47 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_48 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h30 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_48 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_48 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_48 <= btb_510;
      end else begin
        btb_48 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_49 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h31 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_49 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_49 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_49 <= btb_510;
      end else begin
        btb_49 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_50 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h32 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_50 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_50 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_50 <= btb_510;
      end else begin
        btb_50 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_51 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h33 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_51 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_51 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_51 <= btb_510;
      end else begin
        btb_51 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_52 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h34 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_52 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_52 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_52 <= btb_510;
      end else begin
        btb_52 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_53 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h35 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_53 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_53 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_53 <= btb_510;
      end else begin
        btb_53 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_54 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h36 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_54 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_54 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_54 <= btb_510;
      end else begin
        btb_54 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_55 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h37 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_55 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_55 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_55 <= btb_510;
      end else begin
        btb_55 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_56 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h38 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_56 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_56 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_56 <= btb_510;
      end else begin
        btb_56 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_57 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h39 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_57 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_57 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_57 <= btb_510;
      end else begin
        btb_57 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_58 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h3a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_58 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_58 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_58 <= btb_510;
      end else begin
        btb_58 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_59 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h3b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_59 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_59 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_59 <= btb_510;
      end else begin
        btb_59 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_60 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h3c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_60 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_60 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_60 <= btb_510;
      end else begin
        btb_60 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_61 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h3d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_61 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_61 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_61 <= btb_510;
      end else begin
        btb_61 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_62 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h3e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_62 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_62 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_62 <= btb_510;
      end else begin
        btb_62 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_63 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h3f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_63 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_63 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_63 <= btb_510;
      end else begin
        btb_63 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_64 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h40 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_64 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_64 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_64 <= btb_510;
      end else begin
        btb_64 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_65 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h41 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_65 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_65 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_65 <= btb_510;
      end else begin
        btb_65 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_66 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h42 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_66 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_66 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_66 <= btb_510;
      end else begin
        btb_66 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_67 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h43 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_67 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_67 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_67 <= btb_510;
      end else begin
        btb_67 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_68 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h44 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_68 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_68 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_68 <= btb_510;
      end else begin
        btb_68 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_69 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h45 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_69 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_69 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_69 <= btb_510;
      end else begin
        btb_69 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_70 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h46 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_70 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_70 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_70 <= btb_510;
      end else begin
        btb_70 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_71 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h47 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_71 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_71 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_71 <= btb_510;
      end else begin
        btb_71 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_72 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h48 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_72 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_72 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_72 <= btb_510;
      end else begin
        btb_72 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_73 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h49 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_73 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_73 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_73 <= btb_510;
      end else begin
        btb_73 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_74 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h4a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_74 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_74 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_74 <= btb_510;
      end else begin
        btb_74 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_75 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h4b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_75 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_75 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_75 <= btb_510;
      end else begin
        btb_75 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_76 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h4c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_76 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_76 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_76 <= btb_510;
      end else begin
        btb_76 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_77 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h4d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_77 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_77 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_77 <= btb_510;
      end else begin
        btb_77 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_78 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h4e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_78 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_78 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_78 <= btb_510;
      end else begin
        btb_78 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_79 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h4f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_79 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_79 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_79 <= btb_510;
      end else begin
        btb_79 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_80 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h50 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_80 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_80 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_80 <= btb_510;
      end else begin
        btb_80 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_81 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h51 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_81 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_81 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_81 <= btb_510;
      end else begin
        btb_81 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_82 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h52 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_82 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_82 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_82 <= btb_510;
      end else begin
        btb_82 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_83 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h53 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_83 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_83 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_83 <= btb_510;
      end else begin
        btb_83 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_84 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h54 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_84 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_84 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_84 <= btb_510;
      end else begin
        btb_84 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_85 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h55 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_85 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_85 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_85 <= btb_510;
      end else begin
        btb_85 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_86 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h56 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_86 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_86 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_86 <= btb_510;
      end else begin
        btb_86 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_87 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h57 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_87 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_87 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_87 <= btb_510;
      end else begin
        btb_87 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_88 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h58 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_88 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_88 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_88 <= btb_510;
      end else begin
        btb_88 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_89 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h59 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_89 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_89 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_89 <= btb_510;
      end else begin
        btb_89 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_90 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h5a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_90 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_90 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_90 <= btb_510;
      end else begin
        btb_90 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_91 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h5b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_91 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_91 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_91 <= btb_510;
      end else begin
        btb_91 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_92 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h5c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_92 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_92 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_92 <= btb_510;
      end else begin
        btb_92 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_93 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h5d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_93 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_93 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_93 <= btb_510;
      end else begin
        btb_93 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_94 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h5e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_94 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_94 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_94 <= btb_510;
      end else begin
        btb_94 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_95 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h5f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_95 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_95 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_95 <= btb_510;
      end else begin
        btb_95 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_96 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h60 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_96 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_96 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_96 <= btb_510;
      end else begin
        btb_96 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_97 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h61 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_97 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_97 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_97 <= btb_510;
      end else begin
        btb_97 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_98 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h62 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_98 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_98 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_98 <= btb_510;
      end else begin
        btb_98 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_99 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h63 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_99 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_99 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_99 <= btb_510;
      end else begin
        btb_99 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_100 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h64 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_100 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_100 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_100 <= btb_510;
      end else begin
        btb_100 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_101 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h65 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_101 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_101 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_101 <= btb_510;
      end else begin
        btb_101 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_102 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h66 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_102 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_102 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_102 <= btb_510;
      end else begin
        btb_102 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_103 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h67 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_103 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_103 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_103 <= btb_510;
      end else begin
        btb_103 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_104 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h68 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_104 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_104 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_104 <= btb_510;
      end else begin
        btb_104 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_105 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h69 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_105 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_105 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_105 <= btb_510;
      end else begin
        btb_105 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_106 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h6a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_106 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_106 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_106 <= btb_510;
      end else begin
        btb_106 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_107 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h6b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_107 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_107 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_107 <= btb_510;
      end else begin
        btb_107 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_108 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h6c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_108 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_108 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_108 <= btb_510;
      end else begin
        btb_108 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_109 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h6d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_109 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_109 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_109 <= btb_510;
      end else begin
        btb_109 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_110 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h6e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_110 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_110 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_110 <= btb_510;
      end else begin
        btb_110 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_111 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h6f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_111 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_111 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_111 <= btb_510;
      end else begin
        btb_111 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_112 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h70 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_112 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_112 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_112 <= btb_510;
      end else begin
        btb_112 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_113 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h71 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_113 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_113 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_113 <= btb_510;
      end else begin
        btb_113 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_114 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h72 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_114 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_114 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_114 <= btb_510;
      end else begin
        btb_114 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_115 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h73 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_115 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_115 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_115 <= btb_510;
      end else begin
        btb_115 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_116 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h74 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_116 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_116 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_116 <= btb_510;
      end else begin
        btb_116 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_117 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h75 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_117 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_117 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_117 <= btb_510;
      end else begin
        btb_117 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_118 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h76 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_118 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_118 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_118 <= btb_510;
      end else begin
        btb_118 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_119 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h77 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_119 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_119 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_119 <= btb_510;
      end else begin
        btb_119 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_120 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h78 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_120 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_120 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_120 <= btb_510;
      end else begin
        btb_120 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_121 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h79 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_121 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_121 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_121 <= btb_510;
      end else begin
        btb_121 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_122 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h7a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_122 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_122 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_122 <= btb_510;
      end else begin
        btb_122 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_123 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h7b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_123 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_123 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_123 <= btb_510;
      end else begin
        btb_123 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_124 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h7c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_124 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_124 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_124 <= btb_510;
      end else begin
        btb_124 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_125 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h7d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_125 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_125 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_125 <= btb_510;
      end else begin
        btb_125 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_126 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h7e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_126 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_126 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_126 <= btb_510;
      end else begin
        btb_126 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_127 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h7f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_127 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_127 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_127 <= btb_510;
      end else begin
        btb_127 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_128 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h80 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_128 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_128 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_128 <= btb_510;
      end else begin
        btb_128 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_129 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h81 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_129 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_129 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_129 <= btb_510;
      end else begin
        btb_129 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_130 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h82 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_130 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_130 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_130 <= btb_510;
      end else begin
        btb_130 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_131 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h83 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_131 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_131 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_131 <= btb_510;
      end else begin
        btb_131 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_132 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h84 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_132 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_132 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_132 <= btb_510;
      end else begin
        btb_132 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_133 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h85 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_133 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_133 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_133 <= btb_510;
      end else begin
        btb_133 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_134 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h86 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_134 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_134 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_134 <= btb_510;
      end else begin
        btb_134 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_135 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h87 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_135 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_135 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_135 <= btb_510;
      end else begin
        btb_135 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_136 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h88 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_136 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_136 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_136 <= btb_510;
      end else begin
        btb_136 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_137 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h89 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_137 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_137 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_137 <= btb_510;
      end else begin
        btb_137 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_138 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h8a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_138 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_138 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_138 <= btb_510;
      end else begin
        btb_138 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_139 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h8b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_139 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_139 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_139 <= btb_510;
      end else begin
        btb_139 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_140 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h8c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_140 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_140 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_140 <= btb_510;
      end else begin
        btb_140 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_141 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h8d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_141 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_141 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_141 <= btb_510;
      end else begin
        btb_141 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_142 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h8e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_142 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_142 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_142 <= btb_510;
      end else begin
        btb_142 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_143 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h8f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_143 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_143 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_143 <= btb_510;
      end else begin
        btb_143 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_144 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h90 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_144 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_144 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_144 <= btb_510;
      end else begin
        btb_144 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_145 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h91 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_145 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_145 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_145 <= btb_510;
      end else begin
        btb_145 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_146 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h92 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_146 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_146 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_146 <= btb_510;
      end else begin
        btb_146 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_147 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h93 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_147 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_147 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_147 <= btb_510;
      end else begin
        btb_147 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_148 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h94 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_148 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_148 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_148 <= btb_510;
      end else begin
        btb_148 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_149 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h95 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_149 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_149 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_149 <= btb_510;
      end else begin
        btb_149 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_150 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h96 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_150 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_150 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_150 <= btb_510;
      end else begin
        btb_150 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_151 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h97 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_151 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_151 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_151 <= btb_510;
      end else begin
        btb_151 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_152 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h98 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_152 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_152 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_152 <= btb_510;
      end else begin
        btb_152 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_153 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h99 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_153 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_153 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_153 <= btb_510;
      end else begin
        btb_153 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_154 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h9a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_154 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_154 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_154 <= btb_510;
      end else begin
        btb_154 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_155 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h9b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_155 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_155 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_155 <= btb_510;
      end else begin
        btb_155 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_156 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h9c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_156 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_156 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_156 <= btb_510;
      end else begin
        btb_156 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_157 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h9d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_157 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_157 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_157 <= btb_510;
      end else begin
        btb_157 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_158 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h9e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_158 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_158 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_158 <= btb_510;
      end else begin
        btb_158 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_159 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h9f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_159 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_159 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_159 <= btb_510;
      end else begin
        btb_159 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_160 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_160 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_160 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_160 <= btb_510;
      end else begin
        btb_160 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_161 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_161 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_161 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_161 <= btb_510;
      end else begin
        btb_161 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_162 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_162 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_162 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_162 <= btb_510;
      end else begin
        btb_162 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_163 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_163 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_163 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_163 <= btb_510;
      end else begin
        btb_163 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_164 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_164 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_164 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_164 <= btb_510;
      end else begin
        btb_164 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_165 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_165 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_165 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_165 <= btb_510;
      end else begin
        btb_165 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_166 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_166 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_166 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_166 <= btb_510;
      end else begin
        btb_166 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_167 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_167 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_167 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_167 <= btb_510;
      end else begin
        btb_167 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_168 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_168 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_168 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_168 <= btb_510;
      end else begin
        btb_168 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_169 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'ha9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_169 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_169 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_169 <= btb_510;
      end else begin
        btb_169 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_170 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'haa == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_170 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_170 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_170 <= btb_510;
      end else begin
        btb_170 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_171 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hab == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_171 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_171 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_171 <= btb_510;
      end else begin
        btb_171 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_172 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hac == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_172 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_172 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_172 <= btb_510;
      end else begin
        btb_172 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_173 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'had == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_173 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_173 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_173 <= btb_510;
      end else begin
        btb_173 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_174 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hae == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_174 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_174 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_174 <= btb_510;
      end else begin
        btb_174 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_175 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'haf == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_175 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_175 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_175 <= btb_510;
      end else begin
        btb_175 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_176 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_176 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_176 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_176 <= btb_510;
      end else begin
        btb_176 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_177 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_177 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_177 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_177 <= btb_510;
      end else begin
        btb_177 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_178 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_178 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_178 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_178 <= btb_510;
      end else begin
        btb_178 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_179 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_179 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_179 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_179 <= btb_510;
      end else begin
        btb_179 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_180 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_180 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_180 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_180 <= btb_510;
      end else begin
        btb_180 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_181 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_181 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_181 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_181 <= btb_510;
      end else begin
        btb_181 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_182 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_182 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_182 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_182 <= btb_510;
      end else begin
        btb_182 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_183 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_183 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_183 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_183 <= btb_510;
      end else begin
        btb_183 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_184 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_184 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_184 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_184 <= btb_510;
      end else begin
        btb_184 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_185 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hb9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_185 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_185 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_185 <= btb_510;
      end else begin
        btb_185 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_186 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hba == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_186 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_186 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_186 <= btb_510;
      end else begin
        btb_186 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_187 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hbb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_187 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_187 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_187 <= btb_510;
      end else begin
        btb_187 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_188 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hbc == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_188 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_188 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_188 <= btb_510;
      end else begin
        btb_188 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_189 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hbd == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_189 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_189 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_189 <= btb_510;
      end else begin
        btb_189 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_190 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hbe == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_190 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_190 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_190 <= btb_510;
      end else begin
        btb_190 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_191 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hbf == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_191 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_191 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_191 <= btb_510;
      end else begin
        btb_191 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_192 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_192 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_192 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_192 <= btb_510;
      end else begin
        btb_192 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_193 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_193 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_193 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_193 <= btb_510;
      end else begin
        btb_193 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_194 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_194 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_194 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_194 <= btb_510;
      end else begin
        btb_194 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_195 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_195 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_195 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_195 <= btb_510;
      end else begin
        btb_195 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_196 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_196 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_196 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_196 <= btb_510;
      end else begin
        btb_196 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_197 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_197 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_197 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_197 <= btb_510;
      end else begin
        btb_197 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_198 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_198 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_198 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_198 <= btb_510;
      end else begin
        btb_198 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_199 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_199 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_199 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_199 <= btb_510;
      end else begin
        btb_199 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_200 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_200 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_200 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_200 <= btb_510;
      end else begin
        btb_200 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_201 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hc9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_201 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_201 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_201 <= btb_510;
      end else begin
        btb_201 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_202 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hca == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_202 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_202 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_202 <= btb_510;
      end else begin
        btb_202 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_203 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hcb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_203 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_203 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_203 <= btb_510;
      end else begin
        btb_203 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_204 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hcc == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_204 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_204 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_204 <= btb_510;
      end else begin
        btb_204 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_205 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hcd == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_205 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_205 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_205 <= btb_510;
      end else begin
        btb_205 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_206 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hce == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_206 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_206 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_206 <= btb_510;
      end else begin
        btb_206 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_207 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hcf == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_207 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_207 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_207 <= btb_510;
      end else begin
        btb_207 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_208 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_208 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_208 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_208 <= btb_510;
      end else begin
        btb_208 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_209 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_209 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_209 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_209 <= btb_510;
      end else begin
        btb_209 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_210 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_210 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_210 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_210 <= btb_510;
      end else begin
        btb_210 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_211 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_211 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_211 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_211 <= btb_510;
      end else begin
        btb_211 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_212 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_212 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_212 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_212 <= btb_510;
      end else begin
        btb_212 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_213 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_213 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_213 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_213 <= btb_510;
      end else begin
        btb_213 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_214 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_214 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_214 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_214 <= btb_510;
      end else begin
        btb_214 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_215 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_215 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_215 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_215 <= btb_510;
      end else begin
        btb_215 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_216 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_216 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_216 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_216 <= btb_510;
      end else begin
        btb_216 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_217 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hd9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_217 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_217 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_217 <= btb_510;
      end else begin
        btb_217 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_218 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hda == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_218 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_218 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_218 <= btb_510;
      end else begin
        btb_218 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_219 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hdb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_219 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_219 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_219 <= btb_510;
      end else begin
        btb_219 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_220 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hdc == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_220 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_220 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_220 <= btb_510;
      end else begin
        btb_220 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_221 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hdd == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_221 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_221 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_221 <= btb_510;
      end else begin
        btb_221 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_222 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hde == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_222 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_222 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_222 <= btb_510;
      end else begin
        btb_222 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_223 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hdf == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_223 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_223 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_223 <= btb_510;
      end else begin
        btb_223 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_224 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_224 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_224 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_224 <= btb_510;
      end else begin
        btb_224 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_225 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_225 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_225 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_225 <= btb_510;
      end else begin
        btb_225 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_226 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_226 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_226 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_226 <= btb_510;
      end else begin
        btb_226 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_227 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_227 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_227 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_227 <= btb_510;
      end else begin
        btb_227 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_228 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_228 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_228 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_228 <= btb_510;
      end else begin
        btb_228 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_229 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_229 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_229 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_229 <= btb_510;
      end else begin
        btb_229 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_230 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_230 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_230 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_230 <= btb_510;
      end else begin
        btb_230 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_231 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_231 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_231 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_231 <= btb_510;
      end else begin
        btb_231 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_232 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_232 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_232 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_232 <= btb_510;
      end else begin
        btb_232 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_233 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'he9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_233 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_233 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_233 <= btb_510;
      end else begin
        btb_233 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_234 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hea == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_234 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_234 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_234 <= btb_510;
      end else begin
        btb_234 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_235 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'heb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_235 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_235 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_235 <= btb_510;
      end else begin
        btb_235 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_236 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hec == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_236 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_236 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_236 <= btb_510;
      end else begin
        btb_236 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_237 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hed == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_237 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_237 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_237 <= btb_510;
      end else begin
        btb_237 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_238 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hee == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_238 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_238 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_238 <= btb_510;
      end else begin
        btb_238 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_239 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hef == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_239 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_239 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_239 <= btb_510;
      end else begin
        btb_239 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_240 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_240 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_240 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_240 <= btb_510;
      end else begin
        btb_240 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_241 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_241 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_241 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_241 <= btb_510;
      end else begin
        btb_241 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_242 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_242 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_242 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_242 <= btb_510;
      end else begin
        btb_242 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_243 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_243 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_243 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_243 <= btb_510;
      end else begin
        btb_243 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_244 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_244 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_244 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_244 <= btb_510;
      end else begin
        btb_244 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_245 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_245 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_245 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_245 <= btb_510;
      end else begin
        btb_245 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_246 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_246 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_246 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_246 <= btb_510;
      end else begin
        btb_246 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_247 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_247 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_247 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_247 <= btb_510;
      end else begin
        btb_247 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_248 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_248 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_248 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_248 <= btb_510;
      end else begin
        btb_248 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_249 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hf9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_249 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_249 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_249 <= btb_510;
      end else begin
        btb_249 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_250 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hfa == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_250 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_250 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_250 <= btb_510;
      end else begin
        btb_250 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_251 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hfb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_251 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_251 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_251 <= btb_510;
      end else begin
        btb_251 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_252 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hfc == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_252 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_252 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_252 <= btb_510;
      end else begin
        btb_252 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_253 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hfd == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_253 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_253 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_253 <= btb_510;
      end else begin
        btb_253 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_254 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hfe == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_254 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_254 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_254 <= btb_510;
      end else begin
        btb_254 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_255 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'hff == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_255 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_255 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_255 <= btb_510;
      end else begin
        btb_255 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_256 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h100 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_256 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_256 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_256 <= btb_510;
      end else begin
        btb_256 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_257 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h101 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_257 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_257 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_257 <= btb_510;
      end else begin
        btb_257 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_258 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h102 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_258 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_258 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_258 <= btb_510;
      end else begin
        btb_258 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_259 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h103 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_259 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_259 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_259 <= btb_510;
      end else begin
        btb_259 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_260 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h104 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_260 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_260 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_260 <= btb_510;
      end else begin
        btb_260 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_261 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h105 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_261 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_261 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_261 <= btb_510;
      end else begin
        btb_261 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_262 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h106 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_262 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_262 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_262 <= btb_510;
      end else begin
        btb_262 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_263 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h107 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_263 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_263 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_263 <= btb_510;
      end else begin
        btb_263 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_264 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h108 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_264 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_264 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_264 <= btb_510;
      end else begin
        btb_264 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_265 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h109 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_265 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_265 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_265 <= btb_510;
      end else begin
        btb_265 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_266 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h10a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_266 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_266 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_266 <= btb_510;
      end else begin
        btb_266 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_267 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h10b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_267 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_267 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_267 <= btb_510;
      end else begin
        btb_267 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_268 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h10c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_268 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_268 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_268 <= btb_510;
      end else begin
        btb_268 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_269 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h10d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_269 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_269 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_269 <= btb_510;
      end else begin
        btb_269 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_270 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h10e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_270 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_270 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_270 <= btb_510;
      end else begin
        btb_270 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_271 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h10f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_271 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_271 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_271 <= btb_510;
      end else begin
        btb_271 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_272 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h110 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_272 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_272 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_272 <= btb_510;
      end else begin
        btb_272 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_273 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h111 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_273 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_273 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_273 <= btb_510;
      end else begin
        btb_273 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_274 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h112 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_274 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_274 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_274 <= btb_510;
      end else begin
        btb_274 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_275 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h113 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_275 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_275 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_275 <= btb_510;
      end else begin
        btb_275 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_276 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h114 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_276 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_276 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_276 <= btb_510;
      end else begin
        btb_276 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_277 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h115 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_277 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_277 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_277 <= btb_510;
      end else begin
        btb_277 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_278 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h116 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_278 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_278 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_278 <= btb_510;
      end else begin
        btb_278 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_279 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h117 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_279 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_279 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_279 <= btb_510;
      end else begin
        btb_279 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_280 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h118 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_280 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_280 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_280 <= btb_510;
      end else begin
        btb_280 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_281 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h119 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_281 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_281 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_281 <= btb_510;
      end else begin
        btb_281 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_282 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h11a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_282 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_282 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_282 <= btb_510;
      end else begin
        btb_282 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_283 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h11b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_283 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_283 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_283 <= btb_510;
      end else begin
        btb_283 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_284 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h11c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_284 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_284 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_284 <= btb_510;
      end else begin
        btb_284 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_285 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h11d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_285 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_285 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_285 <= btb_510;
      end else begin
        btb_285 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_286 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h11e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_286 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_286 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_286 <= btb_510;
      end else begin
        btb_286 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_287 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h11f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_287 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_287 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_287 <= btb_510;
      end else begin
        btb_287 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_288 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h120 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_288 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_288 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_288 <= btb_510;
      end else begin
        btb_288 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_289 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h121 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_289 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_289 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_289 <= btb_510;
      end else begin
        btb_289 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_290 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h122 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_290 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_290 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_290 <= btb_510;
      end else begin
        btb_290 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_291 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h123 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_291 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_291 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_291 <= btb_510;
      end else begin
        btb_291 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_292 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h124 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_292 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_292 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_292 <= btb_510;
      end else begin
        btb_292 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_293 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h125 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_293 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_293 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_293 <= btb_510;
      end else begin
        btb_293 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_294 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h126 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_294 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_294 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_294 <= btb_510;
      end else begin
        btb_294 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_295 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h127 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_295 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_295 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_295 <= btb_510;
      end else begin
        btb_295 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_296 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h128 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_296 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_296 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_296 <= btb_510;
      end else begin
        btb_296 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_297 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h129 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_297 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_297 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_297 <= btb_510;
      end else begin
        btb_297 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_298 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h12a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_298 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_298 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_298 <= btb_510;
      end else begin
        btb_298 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_299 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h12b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_299 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_299 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_299 <= btb_510;
      end else begin
        btb_299 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_300 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h12c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_300 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_300 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_300 <= btb_510;
      end else begin
        btb_300 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_301 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h12d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_301 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_301 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_301 <= btb_510;
      end else begin
        btb_301 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_302 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h12e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_302 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_302 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_302 <= btb_510;
      end else begin
        btb_302 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_303 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h12f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_303 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_303 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_303 <= btb_510;
      end else begin
        btb_303 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_304 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h130 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_304 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_304 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_304 <= btb_510;
      end else begin
        btb_304 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_305 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h131 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_305 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_305 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_305 <= btb_510;
      end else begin
        btb_305 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_306 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h132 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_306 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_306 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_306 <= btb_510;
      end else begin
        btb_306 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_307 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h133 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_307 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_307 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_307 <= btb_510;
      end else begin
        btb_307 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_308 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h134 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_308 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_308 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_308 <= btb_510;
      end else begin
        btb_308 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_309 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h135 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_309 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_309 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_309 <= btb_510;
      end else begin
        btb_309 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_310 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h136 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_310 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_310 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_310 <= btb_510;
      end else begin
        btb_310 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_311 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h137 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_311 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_311 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_311 <= btb_510;
      end else begin
        btb_311 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_312 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h138 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_312 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_312 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_312 <= btb_510;
      end else begin
        btb_312 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_313 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h139 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_313 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_313 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_313 <= btb_510;
      end else begin
        btb_313 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_314 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h13a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_314 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_314 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_314 <= btb_510;
      end else begin
        btb_314 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_315 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h13b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_315 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_315 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_315 <= btb_510;
      end else begin
        btb_315 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_316 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h13c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_316 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_316 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_316 <= btb_510;
      end else begin
        btb_316 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_317 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h13d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_317 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_317 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_317 <= btb_510;
      end else begin
        btb_317 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_318 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h13e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_318 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_318 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_318 <= btb_510;
      end else begin
        btb_318 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_319 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h13f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_319 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_319 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_319 <= btb_510;
      end else begin
        btb_319 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_320 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h140 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_320 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_320 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_320 <= btb_510;
      end else begin
        btb_320 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_321 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h141 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_321 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_321 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_321 <= btb_510;
      end else begin
        btb_321 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_322 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h142 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_322 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_322 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_322 <= btb_510;
      end else begin
        btb_322 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_323 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h143 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_323 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_323 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_323 <= btb_510;
      end else begin
        btb_323 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_324 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h144 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_324 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_324 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_324 <= btb_510;
      end else begin
        btb_324 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_325 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h145 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_325 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_325 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_325 <= btb_510;
      end else begin
        btb_325 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_326 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h146 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_326 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_326 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_326 <= btb_510;
      end else begin
        btb_326 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_327 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h147 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_327 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_327 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_327 <= btb_510;
      end else begin
        btb_327 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_328 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h148 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_328 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_328 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_328 <= btb_510;
      end else begin
        btb_328 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_329 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h149 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_329 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_329 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_329 <= btb_510;
      end else begin
        btb_329 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_330 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h14a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_330 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_330 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_330 <= btb_510;
      end else begin
        btb_330 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_331 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h14b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_331 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_331 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_331 <= btb_510;
      end else begin
        btb_331 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_332 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h14c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_332 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_332 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_332 <= btb_510;
      end else begin
        btb_332 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_333 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h14d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_333 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_333 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_333 <= btb_510;
      end else begin
        btb_333 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_334 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h14e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_334 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_334 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_334 <= btb_510;
      end else begin
        btb_334 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_335 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h14f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_335 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_335 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_335 <= btb_510;
      end else begin
        btb_335 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_336 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h150 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_336 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_336 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_336 <= btb_510;
      end else begin
        btb_336 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_337 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h151 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_337 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_337 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_337 <= btb_510;
      end else begin
        btb_337 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_338 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h152 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_338 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_338 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_338 <= btb_510;
      end else begin
        btb_338 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_339 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h153 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_339 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_339 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_339 <= btb_510;
      end else begin
        btb_339 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_340 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h154 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_340 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_340 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_340 <= btb_510;
      end else begin
        btb_340 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_341 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h155 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_341 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_341 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_341 <= btb_510;
      end else begin
        btb_341 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_342 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h156 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_342 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_342 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_342 <= btb_510;
      end else begin
        btb_342 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_343 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h157 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_343 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_343 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_343 <= btb_510;
      end else begin
        btb_343 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_344 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h158 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_344 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_344 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_344 <= btb_510;
      end else begin
        btb_344 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_345 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h159 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_345 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_345 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_345 <= btb_510;
      end else begin
        btb_345 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_346 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h15a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_346 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_346 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_346 <= btb_510;
      end else begin
        btb_346 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_347 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h15b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_347 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_347 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_347 <= btb_510;
      end else begin
        btb_347 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_348 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h15c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_348 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_348 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_348 <= btb_510;
      end else begin
        btb_348 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_349 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h15d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_349 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_349 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_349 <= btb_510;
      end else begin
        btb_349 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_350 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h15e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_350 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_350 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_350 <= btb_510;
      end else begin
        btb_350 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_351 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h15f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_351 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_351 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_351 <= btb_510;
      end else begin
        btb_351 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_352 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h160 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_352 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_352 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_352 <= btb_510;
      end else begin
        btb_352 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_353 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h161 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_353 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_353 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_353 <= btb_510;
      end else begin
        btb_353 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_354 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h162 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_354 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_354 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_354 <= btb_510;
      end else begin
        btb_354 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_355 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h163 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_355 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_355 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_355 <= btb_510;
      end else begin
        btb_355 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_356 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h164 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_356 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_356 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_356 <= btb_510;
      end else begin
        btb_356 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_357 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h165 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_357 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_357 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_357 <= btb_510;
      end else begin
        btb_357 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_358 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h166 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_358 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_358 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_358 <= btb_510;
      end else begin
        btb_358 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_359 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h167 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_359 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_359 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_359 <= btb_510;
      end else begin
        btb_359 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_360 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h168 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_360 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_360 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_360 <= btb_510;
      end else begin
        btb_360 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_361 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h169 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_361 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_361 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_361 <= btb_510;
      end else begin
        btb_361 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_362 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h16a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_362 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_362 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_362 <= btb_510;
      end else begin
        btb_362 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_363 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h16b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_363 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_363 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_363 <= btb_510;
      end else begin
        btb_363 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_364 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h16c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_364 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_364 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_364 <= btb_510;
      end else begin
        btb_364 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_365 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h16d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_365 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_365 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_365 <= btb_510;
      end else begin
        btb_365 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_366 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h16e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_366 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_366 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_366 <= btb_510;
      end else begin
        btb_366 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_367 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h16f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_367 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_367 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_367 <= btb_510;
      end else begin
        btb_367 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_368 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h170 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_368 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_368 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_368 <= btb_510;
      end else begin
        btb_368 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_369 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h171 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_369 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_369 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_369 <= btb_510;
      end else begin
        btb_369 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_370 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h172 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_370 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_370 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_370 <= btb_510;
      end else begin
        btb_370 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_371 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h173 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_371 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_371 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_371 <= btb_510;
      end else begin
        btb_371 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_372 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h174 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_372 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_372 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_372 <= btb_510;
      end else begin
        btb_372 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_373 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h175 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_373 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_373 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_373 <= btb_510;
      end else begin
        btb_373 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_374 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h176 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_374 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_374 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_374 <= btb_510;
      end else begin
        btb_374 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_375 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h177 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_375 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_375 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_375 <= btb_510;
      end else begin
        btb_375 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_376 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h178 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_376 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_376 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_376 <= btb_510;
      end else begin
        btb_376 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_377 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h179 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_377 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_377 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_377 <= btb_510;
      end else begin
        btb_377 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_378 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h17a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_378 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_378 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_378 <= btb_510;
      end else begin
        btb_378 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_379 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h17b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_379 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_379 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_379 <= btb_510;
      end else begin
        btb_379 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_380 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h17c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_380 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_380 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_380 <= btb_510;
      end else begin
        btb_380 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_381 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h17d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_381 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_381 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_381 <= btb_510;
      end else begin
        btb_381 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_382 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h17e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_382 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_382 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_382 <= btb_510;
      end else begin
        btb_382 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_383 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h17f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_383 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_383 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_383 <= btb_510;
      end else begin
        btb_383 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_384 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h180 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_384 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_384 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_384 <= btb_510;
      end else begin
        btb_384 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_385 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h181 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_385 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_385 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_385 <= btb_510;
      end else begin
        btb_385 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_386 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h182 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_386 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_386 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_386 <= btb_510;
      end else begin
        btb_386 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_387 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h183 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_387 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_387 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_387 <= btb_510;
      end else begin
        btb_387 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_388 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h184 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_388 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_388 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_388 <= btb_510;
      end else begin
        btb_388 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_389 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h185 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_389 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_389 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_389 <= btb_510;
      end else begin
        btb_389 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_390 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h186 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_390 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_390 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_390 <= btb_510;
      end else begin
        btb_390 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_391 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h187 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_391 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_391 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_391 <= btb_510;
      end else begin
        btb_391 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_392 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h188 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_392 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_392 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_392 <= btb_510;
      end else begin
        btb_392 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_393 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h189 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_393 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_393 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_393 <= btb_510;
      end else begin
        btb_393 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_394 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h18a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_394 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_394 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_394 <= btb_510;
      end else begin
        btb_394 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_395 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h18b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_395 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_395 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_395 <= btb_510;
      end else begin
        btb_395 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_396 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h18c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_396 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_396 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_396 <= btb_510;
      end else begin
        btb_396 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_397 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h18d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_397 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_397 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_397 <= btb_510;
      end else begin
        btb_397 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_398 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h18e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_398 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_398 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_398 <= btb_510;
      end else begin
        btb_398 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_399 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h18f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_399 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_399 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_399 <= btb_510;
      end else begin
        btb_399 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_400 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h190 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_400 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_400 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_400 <= btb_510;
      end else begin
        btb_400 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_401 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h191 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_401 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_401 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_401 <= btb_510;
      end else begin
        btb_401 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_402 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h192 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_402 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_402 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_402 <= btb_510;
      end else begin
        btb_402 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_403 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h193 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_403 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_403 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_403 <= btb_510;
      end else begin
        btb_403 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_404 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h194 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_404 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_404 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_404 <= btb_510;
      end else begin
        btb_404 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_405 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h195 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_405 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_405 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_405 <= btb_510;
      end else begin
        btb_405 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_406 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h196 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_406 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_406 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_406 <= btb_510;
      end else begin
        btb_406 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_407 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h197 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_407 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_407 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_407 <= btb_510;
      end else begin
        btb_407 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_408 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h198 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_408 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_408 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_408 <= btb_510;
      end else begin
        btb_408 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_409 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h199 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_409 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_409 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_409 <= btb_510;
      end else begin
        btb_409 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_410 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h19a == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_410 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_410 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_410 <= btb_510;
      end else begin
        btb_410 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_411 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h19b == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_411 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_411 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_411 <= btb_510;
      end else begin
        btb_411 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_412 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h19c == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_412 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_412 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_412 <= btb_510;
      end else begin
        btb_412 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_413 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h19d == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_413 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_413 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_413 <= btb_510;
      end else begin
        btb_413 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_414 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h19e == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_414 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_414 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_414 <= btb_510;
      end else begin
        btb_414 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_415 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h19f == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_415 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_415 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_415 <= btb_510;
      end else begin
        btb_415 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_416 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_416 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_416 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_416 <= btb_510;
      end else begin
        btb_416 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_417 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_417 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_417 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_417 <= btb_510;
      end else begin
        btb_417 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_418 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_418 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_418 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_418 <= btb_510;
      end else begin
        btb_418 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_419 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_419 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_419 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_419 <= btb_510;
      end else begin
        btb_419 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_420 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_420 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_420 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_420 <= btb_510;
      end else begin
        btb_420 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_421 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_421 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_421 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_421 <= btb_510;
      end else begin
        btb_421 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_422 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_422 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_422 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_422 <= btb_510;
      end else begin
        btb_422 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_423 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_423 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_423 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_423 <= btb_510;
      end else begin
        btb_423 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_424 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_424 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_424 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_424 <= btb_510;
      end else begin
        btb_424 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_425 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1a9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_425 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_425 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_425 <= btb_510;
      end else begin
        btb_425 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_426 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1aa == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_426 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_426 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_426 <= btb_510;
      end else begin
        btb_426 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_427 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ab == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_427 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_427 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_427 <= btb_510;
      end else begin
        btb_427 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_428 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ac == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_428 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_428 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_428 <= btb_510;
      end else begin
        btb_428 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_429 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ad == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_429 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_429 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_429 <= btb_510;
      end else begin
        btb_429 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_430 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ae == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_430 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_430 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_430 <= btb_510;
      end else begin
        btb_430 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_431 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1af == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_431 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_431 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_431 <= btb_510;
      end else begin
        btb_431 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_432 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_432 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_432 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_432 <= btb_510;
      end else begin
        btb_432 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_433 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_433 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_433 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_433 <= btb_510;
      end else begin
        btb_433 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_434 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_434 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_434 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_434 <= btb_510;
      end else begin
        btb_434 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_435 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_435 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_435 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_435 <= btb_510;
      end else begin
        btb_435 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_436 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_436 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_436 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_436 <= btb_510;
      end else begin
        btb_436 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_437 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_437 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_437 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_437 <= btb_510;
      end else begin
        btb_437 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_438 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_438 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_438 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_438 <= btb_510;
      end else begin
        btb_438 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_439 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_439 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_439 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_439 <= btb_510;
      end else begin
        btb_439 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_440 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_440 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_440 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_440 <= btb_510;
      end else begin
        btb_440 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_441 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1b9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_441 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_441 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_441 <= btb_510;
      end else begin
        btb_441 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_442 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ba == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_442 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_442 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_442 <= btb_510;
      end else begin
        btb_442 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_443 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1bb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_443 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_443 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_443 <= btb_510;
      end else begin
        btb_443 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_444 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1bc == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_444 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_444 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_444 <= btb_510;
      end else begin
        btb_444 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_445 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1bd == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_445 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_445 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_445 <= btb_510;
      end else begin
        btb_445 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_446 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1be == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_446 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_446 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_446 <= btb_510;
      end else begin
        btb_446 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_447 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1bf == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_447 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_447 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_447 <= btb_510;
      end else begin
        btb_447 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_448 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_448 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_448 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_448 <= btb_510;
      end else begin
        btb_448 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_449 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_449 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_449 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_449 <= btb_510;
      end else begin
        btb_449 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_450 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_450 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_450 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_450 <= btb_510;
      end else begin
        btb_450 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_451 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_451 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_451 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_451 <= btb_510;
      end else begin
        btb_451 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_452 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_452 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_452 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_452 <= btb_510;
      end else begin
        btb_452 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_453 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_453 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_453 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_453 <= btb_510;
      end else begin
        btb_453 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_454 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_454 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_454 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_454 <= btb_510;
      end else begin
        btb_454 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_455 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_455 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_455 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_455 <= btb_510;
      end else begin
        btb_455 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_456 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_456 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_456 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_456 <= btb_510;
      end else begin
        btb_456 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_457 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1c9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_457 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_457 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_457 <= btb_510;
      end else begin
        btb_457 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_458 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ca == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_458 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_458 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_458 <= btb_510;
      end else begin
        btb_458 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_459 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1cb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_459 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_459 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_459 <= btb_510;
      end else begin
        btb_459 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_460 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1cc == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_460 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_460 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_460 <= btb_510;
      end else begin
        btb_460 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_461 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1cd == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_461 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_461 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_461 <= btb_510;
      end else begin
        btb_461 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_462 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ce == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_462 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_462 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_462 <= btb_510;
      end else begin
        btb_462 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_463 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1cf == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_463 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_463 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_463 <= btb_510;
      end else begin
        btb_463 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_464 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_464 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_464 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_464 <= btb_510;
      end else begin
        btb_464 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_465 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_465 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_465 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_465 <= btb_510;
      end else begin
        btb_465 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_466 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_466 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_466 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_466 <= btb_510;
      end else begin
        btb_466 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_467 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_467 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_467 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_467 <= btb_510;
      end else begin
        btb_467 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_468 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_468 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_468 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_468 <= btb_510;
      end else begin
        btb_468 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_469 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_469 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_469 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_469 <= btb_510;
      end else begin
        btb_469 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_470 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_470 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_470 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_470 <= btb_510;
      end else begin
        btb_470 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_471 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_471 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_471 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_471 <= btb_510;
      end else begin
        btb_471 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_472 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_472 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_472 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_472 <= btb_510;
      end else begin
        btb_472 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_473 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1d9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_473 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_473 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_473 <= btb_510;
      end else begin
        btb_473 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_474 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1da == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_474 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_474 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_474 <= btb_510;
      end else begin
        btb_474 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_475 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1db == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_475 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_475 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_475 <= btb_510;
      end else begin
        btb_475 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_476 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1dc == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_476 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_476 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_476 <= btb_510;
      end else begin
        btb_476 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_477 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1dd == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_477 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_477 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_477 <= btb_510;
      end else begin
        btb_477 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_478 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1de == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_478 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_478 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_478 <= btb_510;
      end else begin
        btb_478 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_479 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1df == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_479 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_479 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_479 <= btb_510;
      end else begin
        btb_479 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_480 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_480 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_480 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_480 <= btb_510;
      end else begin
        btb_480 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_481 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_481 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_481 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_481 <= btb_510;
      end else begin
        btb_481 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_482 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_482 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_482 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_482 <= btb_510;
      end else begin
        btb_482 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_483 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_483 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_483 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_483 <= btb_510;
      end else begin
        btb_483 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_484 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_484 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_484 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_484 <= btb_510;
      end else begin
        btb_484 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_485 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_485 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_485 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_485 <= btb_510;
      end else begin
        btb_485 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_486 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_486 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_486 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_486 <= btb_510;
      end else begin
        btb_486 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_487 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_487 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_487 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_487 <= btb_510;
      end else begin
        btb_487 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_488 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_488 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_488 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_488 <= btb_510;
      end else begin
        btb_488 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_489 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1e9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_489 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_489 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_489 <= btb_510;
      end else begin
        btb_489 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_490 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ea == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_490 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_490 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_490 <= btb_510;
      end else begin
        btb_490 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_491 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1eb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_491 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_491 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_491 <= btb_510;
      end else begin
        btb_491 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_492 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ec == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_492 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_492 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_492 <= btb_510;
      end else begin
        btb_492 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_493 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ed == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_493 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_493 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_493 <= btb_510;
      end else begin
        btb_493 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_494 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ee == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_494 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_494 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_494 <= btb_510;
      end else begin
        btb_494 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_495 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ef == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_495 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_495 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_495 <= btb_510;
      end else begin
        btb_495 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_496 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f0 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_496 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_496 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_496 <= btb_510;
      end else begin
        btb_496 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_497 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f1 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_497 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_497 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_497 <= btb_510;
      end else begin
        btb_497 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_498 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f2 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_498 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_498 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_498 <= btb_510;
      end else begin
        btb_498 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_499 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f3 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_499 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_499 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_499 <= btb_510;
      end else begin
        btb_499 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_500 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f4 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_500 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_500 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_500 <= btb_510;
      end else begin
        btb_500 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_501 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f5 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_501 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_501 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_501 <= btb_510;
      end else begin
        btb_501 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_502 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f6 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_502 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_502 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_502 <= btb_510;
      end else begin
        btb_502 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_503 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f7 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_503 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_503 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_503 <= btb_510;
      end else begin
        btb_503 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_504 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f8 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_504 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_504 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_504 <= btb_510;
      end else begin
        btb_504 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_505 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1f9 == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_505 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_505 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_505 <= btb_510;
      end else begin
        btb_505 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_506 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1fa == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_506 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_506 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_506 <= btb_510;
      end else begin
        btb_506 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_507 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1fb == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_507 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_507 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_507 <= btb_510;
      end else begin
        btb_507 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_508 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1fc == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_508 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_508 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_508 <= btb_510;
      end else begin
        btb_508 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_509 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1fd == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_509 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_509 <= btb_511;
      end else if (9'h1fe == io_aw_addr) begin
        btb_509 <= btb_510;
      end else begin
        btb_509 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_510 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1fe == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_510 <= io_in;
      end else if (9'h1ff == io_aw_addr) begin
        btb_510 <= btb_511;
      end else if (!(9'h1fe == io_aw_addr)) begin
        btb_510 <= _GEN_1021;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[ports_lookup_table.scala 83:21]
      btb_511 <= 32'h0; // @[ports_lookup_table.scala 83:{27,27,27,27,27}]
    end else if (9'h1ff == io_aw_addr) begin // @[ports_lookup_table.scala 81:22]
      if (io_write) begin
        btb_511 <= io_in;
      end else if (!(9'h1ff == io_aw_addr)) begin
        if (9'h1fe == io_aw_addr) begin
          btb_511 <= btb_510;
        end else begin
          btb_511 <= _GEN_1021;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  btb_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  btb_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  btb_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  btb_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  btb_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  btb_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  btb_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  btb_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  btb_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  btb_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  btb_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  btb_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  btb_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  btb_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  btb_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  btb_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  btb_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  btb_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  btb_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  btb_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  btb_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  btb_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  btb_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  btb_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  btb_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  btb_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  btb_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  btb_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  btb_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  btb_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  btb_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  btb_31 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  btb_32 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  btb_33 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  btb_34 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  btb_35 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  btb_36 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  btb_37 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  btb_38 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  btb_39 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  btb_40 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  btb_41 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  btb_42 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  btb_43 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  btb_44 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  btb_45 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  btb_46 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  btb_47 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  btb_48 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  btb_49 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  btb_50 = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  btb_51 = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  btb_52 = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  btb_53 = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  btb_54 = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  btb_55 = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  btb_56 = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  btb_57 = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  btb_58 = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  btb_59 = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  btb_60 = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  btb_61 = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  btb_62 = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  btb_63 = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  btb_64 = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  btb_65 = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  btb_66 = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  btb_67 = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  btb_68 = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  btb_69 = _RAND_69[31:0];
  _RAND_70 = {1{`RANDOM}};
  btb_70 = _RAND_70[31:0];
  _RAND_71 = {1{`RANDOM}};
  btb_71 = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  btb_72 = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  btb_73 = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  btb_74 = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  btb_75 = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  btb_76 = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  btb_77 = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  btb_78 = _RAND_78[31:0];
  _RAND_79 = {1{`RANDOM}};
  btb_79 = _RAND_79[31:0];
  _RAND_80 = {1{`RANDOM}};
  btb_80 = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  btb_81 = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  btb_82 = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  btb_83 = _RAND_83[31:0];
  _RAND_84 = {1{`RANDOM}};
  btb_84 = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  btb_85 = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  btb_86 = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  btb_87 = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  btb_88 = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  btb_89 = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  btb_90 = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  btb_91 = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  btb_92 = _RAND_92[31:0];
  _RAND_93 = {1{`RANDOM}};
  btb_93 = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  btb_94 = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  btb_95 = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  btb_96 = _RAND_96[31:0];
  _RAND_97 = {1{`RANDOM}};
  btb_97 = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  btb_98 = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  btb_99 = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  btb_100 = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  btb_101 = _RAND_101[31:0];
  _RAND_102 = {1{`RANDOM}};
  btb_102 = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  btb_103 = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  btb_104 = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  btb_105 = _RAND_105[31:0];
  _RAND_106 = {1{`RANDOM}};
  btb_106 = _RAND_106[31:0];
  _RAND_107 = {1{`RANDOM}};
  btb_107 = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  btb_108 = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  btb_109 = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  btb_110 = _RAND_110[31:0];
  _RAND_111 = {1{`RANDOM}};
  btb_111 = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  btb_112 = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  btb_113 = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  btb_114 = _RAND_114[31:0];
  _RAND_115 = {1{`RANDOM}};
  btb_115 = _RAND_115[31:0];
  _RAND_116 = {1{`RANDOM}};
  btb_116 = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  btb_117 = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  btb_118 = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  btb_119 = _RAND_119[31:0];
  _RAND_120 = {1{`RANDOM}};
  btb_120 = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  btb_121 = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  btb_122 = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  btb_123 = _RAND_123[31:0];
  _RAND_124 = {1{`RANDOM}};
  btb_124 = _RAND_124[31:0];
  _RAND_125 = {1{`RANDOM}};
  btb_125 = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  btb_126 = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  btb_127 = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  btb_128 = _RAND_128[31:0];
  _RAND_129 = {1{`RANDOM}};
  btb_129 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  btb_130 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  btb_131 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  btb_132 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  btb_133 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  btb_134 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  btb_135 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  btb_136 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  btb_137 = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  btb_138 = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  btb_139 = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  btb_140 = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  btb_141 = _RAND_141[31:0];
  _RAND_142 = {1{`RANDOM}};
  btb_142 = _RAND_142[31:0];
  _RAND_143 = {1{`RANDOM}};
  btb_143 = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  btb_144 = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  btb_145 = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  btb_146 = _RAND_146[31:0];
  _RAND_147 = {1{`RANDOM}};
  btb_147 = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  btb_148 = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  btb_149 = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  btb_150 = _RAND_150[31:0];
  _RAND_151 = {1{`RANDOM}};
  btb_151 = _RAND_151[31:0];
  _RAND_152 = {1{`RANDOM}};
  btb_152 = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  btb_153 = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  btb_154 = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  btb_155 = _RAND_155[31:0];
  _RAND_156 = {1{`RANDOM}};
  btb_156 = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  btb_157 = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  btb_158 = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  btb_159 = _RAND_159[31:0];
  _RAND_160 = {1{`RANDOM}};
  btb_160 = _RAND_160[31:0];
  _RAND_161 = {1{`RANDOM}};
  btb_161 = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  btb_162 = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  btb_163 = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  btb_164 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  btb_165 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  btb_166 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  btb_167 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  btb_168 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  btb_169 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  btb_170 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  btb_171 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  btb_172 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  btb_173 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  btb_174 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  btb_175 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  btb_176 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  btb_177 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  btb_178 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  btb_179 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  btb_180 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  btb_181 = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  btb_182 = _RAND_182[31:0];
  _RAND_183 = {1{`RANDOM}};
  btb_183 = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  btb_184 = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  btb_185 = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  btb_186 = _RAND_186[31:0];
  _RAND_187 = {1{`RANDOM}};
  btb_187 = _RAND_187[31:0];
  _RAND_188 = {1{`RANDOM}};
  btb_188 = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  btb_189 = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  btb_190 = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  btb_191 = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  btb_192 = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  btb_193 = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  btb_194 = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  btb_195 = _RAND_195[31:0];
  _RAND_196 = {1{`RANDOM}};
  btb_196 = _RAND_196[31:0];
  _RAND_197 = {1{`RANDOM}};
  btb_197 = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  btb_198 = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  btb_199 = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  btb_200 = _RAND_200[31:0];
  _RAND_201 = {1{`RANDOM}};
  btb_201 = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  btb_202 = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  btb_203 = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  btb_204 = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  btb_205 = _RAND_205[31:0];
  _RAND_206 = {1{`RANDOM}};
  btb_206 = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  btb_207 = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  btb_208 = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  btb_209 = _RAND_209[31:0];
  _RAND_210 = {1{`RANDOM}};
  btb_210 = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  btb_211 = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  btb_212 = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  btb_213 = _RAND_213[31:0];
  _RAND_214 = {1{`RANDOM}};
  btb_214 = _RAND_214[31:0];
  _RAND_215 = {1{`RANDOM}};
  btb_215 = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  btb_216 = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  btb_217 = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  btb_218 = _RAND_218[31:0];
  _RAND_219 = {1{`RANDOM}};
  btb_219 = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  btb_220 = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  btb_221 = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  btb_222 = _RAND_222[31:0];
  _RAND_223 = {1{`RANDOM}};
  btb_223 = _RAND_223[31:0];
  _RAND_224 = {1{`RANDOM}};
  btb_224 = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  btb_225 = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  btb_226 = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  btb_227 = _RAND_227[31:0];
  _RAND_228 = {1{`RANDOM}};
  btb_228 = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  btb_229 = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  btb_230 = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  btb_231 = _RAND_231[31:0];
  _RAND_232 = {1{`RANDOM}};
  btb_232 = _RAND_232[31:0];
  _RAND_233 = {1{`RANDOM}};
  btb_233 = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  btb_234 = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  btb_235 = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  btb_236 = _RAND_236[31:0];
  _RAND_237 = {1{`RANDOM}};
  btb_237 = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  btb_238 = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  btb_239 = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  btb_240 = _RAND_240[31:0];
  _RAND_241 = {1{`RANDOM}};
  btb_241 = _RAND_241[31:0];
  _RAND_242 = {1{`RANDOM}};
  btb_242 = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  btb_243 = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  btb_244 = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  btb_245 = _RAND_245[31:0];
  _RAND_246 = {1{`RANDOM}};
  btb_246 = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  btb_247 = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  btb_248 = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  btb_249 = _RAND_249[31:0];
  _RAND_250 = {1{`RANDOM}};
  btb_250 = _RAND_250[31:0];
  _RAND_251 = {1{`RANDOM}};
  btb_251 = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  btb_252 = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  btb_253 = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  btb_254 = _RAND_254[31:0];
  _RAND_255 = {1{`RANDOM}};
  btb_255 = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  btb_256 = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  btb_257 = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  btb_258 = _RAND_258[31:0];
  _RAND_259 = {1{`RANDOM}};
  btb_259 = _RAND_259[31:0];
  _RAND_260 = {1{`RANDOM}};
  btb_260 = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  btb_261 = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  btb_262 = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  btb_263 = _RAND_263[31:0];
  _RAND_264 = {1{`RANDOM}};
  btb_264 = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  btb_265 = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  btb_266 = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  btb_267 = _RAND_267[31:0];
  _RAND_268 = {1{`RANDOM}};
  btb_268 = _RAND_268[31:0];
  _RAND_269 = {1{`RANDOM}};
  btb_269 = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  btb_270 = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  btb_271 = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  btb_272 = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  btb_273 = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  btb_274 = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  btb_275 = _RAND_275[31:0];
  _RAND_276 = {1{`RANDOM}};
  btb_276 = _RAND_276[31:0];
  _RAND_277 = {1{`RANDOM}};
  btb_277 = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  btb_278 = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  btb_279 = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  btb_280 = _RAND_280[31:0];
  _RAND_281 = {1{`RANDOM}};
  btb_281 = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  btb_282 = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  btb_283 = _RAND_283[31:0];
  _RAND_284 = {1{`RANDOM}};
  btb_284 = _RAND_284[31:0];
  _RAND_285 = {1{`RANDOM}};
  btb_285 = _RAND_285[31:0];
  _RAND_286 = {1{`RANDOM}};
  btb_286 = _RAND_286[31:0];
  _RAND_287 = {1{`RANDOM}};
  btb_287 = _RAND_287[31:0];
  _RAND_288 = {1{`RANDOM}};
  btb_288 = _RAND_288[31:0];
  _RAND_289 = {1{`RANDOM}};
  btb_289 = _RAND_289[31:0];
  _RAND_290 = {1{`RANDOM}};
  btb_290 = _RAND_290[31:0];
  _RAND_291 = {1{`RANDOM}};
  btb_291 = _RAND_291[31:0];
  _RAND_292 = {1{`RANDOM}};
  btb_292 = _RAND_292[31:0];
  _RAND_293 = {1{`RANDOM}};
  btb_293 = _RAND_293[31:0];
  _RAND_294 = {1{`RANDOM}};
  btb_294 = _RAND_294[31:0];
  _RAND_295 = {1{`RANDOM}};
  btb_295 = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  btb_296 = _RAND_296[31:0];
  _RAND_297 = {1{`RANDOM}};
  btb_297 = _RAND_297[31:0];
  _RAND_298 = {1{`RANDOM}};
  btb_298 = _RAND_298[31:0];
  _RAND_299 = {1{`RANDOM}};
  btb_299 = _RAND_299[31:0];
  _RAND_300 = {1{`RANDOM}};
  btb_300 = _RAND_300[31:0];
  _RAND_301 = {1{`RANDOM}};
  btb_301 = _RAND_301[31:0];
  _RAND_302 = {1{`RANDOM}};
  btb_302 = _RAND_302[31:0];
  _RAND_303 = {1{`RANDOM}};
  btb_303 = _RAND_303[31:0];
  _RAND_304 = {1{`RANDOM}};
  btb_304 = _RAND_304[31:0];
  _RAND_305 = {1{`RANDOM}};
  btb_305 = _RAND_305[31:0];
  _RAND_306 = {1{`RANDOM}};
  btb_306 = _RAND_306[31:0];
  _RAND_307 = {1{`RANDOM}};
  btb_307 = _RAND_307[31:0];
  _RAND_308 = {1{`RANDOM}};
  btb_308 = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  btb_309 = _RAND_309[31:0];
  _RAND_310 = {1{`RANDOM}};
  btb_310 = _RAND_310[31:0];
  _RAND_311 = {1{`RANDOM}};
  btb_311 = _RAND_311[31:0];
  _RAND_312 = {1{`RANDOM}};
  btb_312 = _RAND_312[31:0];
  _RAND_313 = {1{`RANDOM}};
  btb_313 = _RAND_313[31:0];
  _RAND_314 = {1{`RANDOM}};
  btb_314 = _RAND_314[31:0];
  _RAND_315 = {1{`RANDOM}};
  btb_315 = _RAND_315[31:0];
  _RAND_316 = {1{`RANDOM}};
  btb_316 = _RAND_316[31:0];
  _RAND_317 = {1{`RANDOM}};
  btb_317 = _RAND_317[31:0];
  _RAND_318 = {1{`RANDOM}};
  btb_318 = _RAND_318[31:0];
  _RAND_319 = {1{`RANDOM}};
  btb_319 = _RAND_319[31:0];
  _RAND_320 = {1{`RANDOM}};
  btb_320 = _RAND_320[31:0];
  _RAND_321 = {1{`RANDOM}};
  btb_321 = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  btb_322 = _RAND_322[31:0];
  _RAND_323 = {1{`RANDOM}};
  btb_323 = _RAND_323[31:0];
  _RAND_324 = {1{`RANDOM}};
  btb_324 = _RAND_324[31:0];
  _RAND_325 = {1{`RANDOM}};
  btb_325 = _RAND_325[31:0];
  _RAND_326 = {1{`RANDOM}};
  btb_326 = _RAND_326[31:0];
  _RAND_327 = {1{`RANDOM}};
  btb_327 = _RAND_327[31:0];
  _RAND_328 = {1{`RANDOM}};
  btb_328 = _RAND_328[31:0];
  _RAND_329 = {1{`RANDOM}};
  btb_329 = _RAND_329[31:0];
  _RAND_330 = {1{`RANDOM}};
  btb_330 = _RAND_330[31:0];
  _RAND_331 = {1{`RANDOM}};
  btb_331 = _RAND_331[31:0];
  _RAND_332 = {1{`RANDOM}};
  btb_332 = _RAND_332[31:0];
  _RAND_333 = {1{`RANDOM}};
  btb_333 = _RAND_333[31:0];
  _RAND_334 = {1{`RANDOM}};
  btb_334 = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  btb_335 = _RAND_335[31:0];
  _RAND_336 = {1{`RANDOM}};
  btb_336 = _RAND_336[31:0];
  _RAND_337 = {1{`RANDOM}};
  btb_337 = _RAND_337[31:0];
  _RAND_338 = {1{`RANDOM}};
  btb_338 = _RAND_338[31:0];
  _RAND_339 = {1{`RANDOM}};
  btb_339 = _RAND_339[31:0];
  _RAND_340 = {1{`RANDOM}};
  btb_340 = _RAND_340[31:0];
  _RAND_341 = {1{`RANDOM}};
  btb_341 = _RAND_341[31:0];
  _RAND_342 = {1{`RANDOM}};
  btb_342 = _RAND_342[31:0];
  _RAND_343 = {1{`RANDOM}};
  btb_343 = _RAND_343[31:0];
  _RAND_344 = {1{`RANDOM}};
  btb_344 = _RAND_344[31:0];
  _RAND_345 = {1{`RANDOM}};
  btb_345 = _RAND_345[31:0];
  _RAND_346 = {1{`RANDOM}};
  btb_346 = _RAND_346[31:0];
  _RAND_347 = {1{`RANDOM}};
  btb_347 = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  btb_348 = _RAND_348[31:0];
  _RAND_349 = {1{`RANDOM}};
  btb_349 = _RAND_349[31:0];
  _RAND_350 = {1{`RANDOM}};
  btb_350 = _RAND_350[31:0];
  _RAND_351 = {1{`RANDOM}};
  btb_351 = _RAND_351[31:0];
  _RAND_352 = {1{`RANDOM}};
  btb_352 = _RAND_352[31:0];
  _RAND_353 = {1{`RANDOM}};
  btb_353 = _RAND_353[31:0];
  _RAND_354 = {1{`RANDOM}};
  btb_354 = _RAND_354[31:0];
  _RAND_355 = {1{`RANDOM}};
  btb_355 = _RAND_355[31:0];
  _RAND_356 = {1{`RANDOM}};
  btb_356 = _RAND_356[31:0];
  _RAND_357 = {1{`RANDOM}};
  btb_357 = _RAND_357[31:0];
  _RAND_358 = {1{`RANDOM}};
  btb_358 = _RAND_358[31:0];
  _RAND_359 = {1{`RANDOM}};
  btb_359 = _RAND_359[31:0];
  _RAND_360 = {1{`RANDOM}};
  btb_360 = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  btb_361 = _RAND_361[31:0];
  _RAND_362 = {1{`RANDOM}};
  btb_362 = _RAND_362[31:0];
  _RAND_363 = {1{`RANDOM}};
  btb_363 = _RAND_363[31:0];
  _RAND_364 = {1{`RANDOM}};
  btb_364 = _RAND_364[31:0];
  _RAND_365 = {1{`RANDOM}};
  btb_365 = _RAND_365[31:0];
  _RAND_366 = {1{`RANDOM}};
  btb_366 = _RAND_366[31:0];
  _RAND_367 = {1{`RANDOM}};
  btb_367 = _RAND_367[31:0];
  _RAND_368 = {1{`RANDOM}};
  btb_368 = _RAND_368[31:0];
  _RAND_369 = {1{`RANDOM}};
  btb_369 = _RAND_369[31:0];
  _RAND_370 = {1{`RANDOM}};
  btb_370 = _RAND_370[31:0];
  _RAND_371 = {1{`RANDOM}};
  btb_371 = _RAND_371[31:0];
  _RAND_372 = {1{`RANDOM}};
  btb_372 = _RAND_372[31:0];
  _RAND_373 = {1{`RANDOM}};
  btb_373 = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  btb_374 = _RAND_374[31:0];
  _RAND_375 = {1{`RANDOM}};
  btb_375 = _RAND_375[31:0];
  _RAND_376 = {1{`RANDOM}};
  btb_376 = _RAND_376[31:0];
  _RAND_377 = {1{`RANDOM}};
  btb_377 = _RAND_377[31:0];
  _RAND_378 = {1{`RANDOM}};
  btb_378 = _RAND_378[31:0];
  _RAND_379 = {1{`RANDOM}};
  btb_379 = _RAND_379[31:0];
  _RAND_380 = {1{`RANDOM}};
  btb_380 = _RAND_380[31:0];
  _RAND_381 = {1{`RANDOM}};
  btb_381 = _RAND_381[31:0];
  _RAND_382 = {1{`RANDOM}};
  btb_382 = _RAND_382[31:0];
  _RAND_383 = {1{`RANDOM}};
  btb_383 = _RAND_383[31:0];
  _RAND_384 = {1{`RANDOM}};
  btb_384 = _RAND_384[31:0];
  _RAND_385 = {1{`RANDOM}};
  btb_385 = _RAND_385[31:0];
  _RAND_386 = {1{`RANDOM}};
  btb_386 = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  btb_387 = _RAND_387[31:0];
  _RAND_388 = {1{`RANDOM}};
  btb_388 = _RAND_388[31:0];
  _RAND_389 = {1{`RANDOM}};
  btb_389 = _RAND_389[31:0];
  _RAND_390 = {1{`RANDOM}};
  btb_390 = _RAND_390[31:0];
  _RAND_391 = {1{`RANDOM}};
  btb_391 = _RAND_391[31:0];
  _RAND_392 = {1{`RANDOM}};
  btb_392 = _RAND_392[31:0];
  _RAND_393 = {1{`RANDOM}};
  btb_393 = _RAND_393[31:0];
  _RAND_394 = {1{`RANDOM}};
  btb_394 = _RAND_394[31:0];
  _RAND_395 = {1{`RANDOM}};
  btb_395 = _RAND_395[31:0];
  _RAND_396 = {1{`RANDOM}};
  btb_396 = _RAND_396[31:0];
  _RAND_397 = {1{`RANDOM}};
  btb_397 = _RAND_397[31:0];
  _RAND_398 = {1{`RANDOM}};
  btb_398 = _RAND_398[31:0];
  _RAND_399 = {1{`RANDOM}};
  btb_399 = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  btb_400 = _RAND_400[31:0];
  _RAND_401 = {1{`RANDOM}};
  btb_401 = _RAND_401[31:0];
  _RAND_402 = {1{`RANDOM}};
  btb_402 = _RAND_402[31:0];
  _RAND_403 = {1{`RANDOM}};
  btb_403 = _RAND_403[31:0];
  _RAND_404 = {1{`RANDOM}};
  btb_404 = _RAND_404[31:0];
  _RAND_405 = {1{`RANDOM}};
  btb_405 = _RAND_405[31:0];
  _RAND_406 = {1{`RANDOM}};
  btb_406 = _RAND_406[31:0];
  _RAND_407 = {1{`RANDOM}};
  btb_407 = _RAND_407[31:0];
  _RAND_408 = {1{`RANDOM}};
  btb_408 = _RAND_408[31:0];
  _RAND_409 = {1{`RANDOM}};
  btb_409 = _RAND_409[31:0];
  _RAND_410 = {1{`RANDOM}};
  btb_410 = _RAND_410[31:0];
  _RAND_411 = {1{`RANDOM}};
  btb_411 = _RAND_411[31:0];
  _RAND_412 = {1{`RANDOM}};
  btb_412 = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  btb_413 = _RAND_413[31:0];
  _RAND_414 = {1{`RANDOM}};
  btb_414 = _RAND_414[31:0];
  _RAND_415 = {1{`RANDOM}};
  btb_415 = _RAND_415[31:0];
  _RAND_416 = {1{`RANDOM}};
  btb_416 = _RAND_416[31:0];
  _RAND_417 = {1{`RANDOM}};
  btb_417 = _RAND_417[31:0];
  _RAND_418 = {1{`RANDOM}};
  btb_418 = _RAND_418[31:0];
  _RAND_419 = {1{`RANDOM}};
  btb_419 = _RAND_419[31:0];
  _RAND_420 = {1{`RANDOM}};
  btb_420 = _RAND_420[31:0];
  _RAND_421 = {1{`RANDOM}};
  btb_421 = _RAND_421[31:0];
  _RAND_422 = {1{`RANDOM}};
  btb_422 = _RAND_422[31:0];
  _RAND_423 = {1{`RANDOM}};
  btb_423 = _RAND_423[31:0];
  _RAND_424 = {1{`RANDOM}};
  btb_424 = _RAND_424[31:0];
  _RAND_425 = {1{`RANDOM}};
  btb_425 = _RAND_425[31:0];
  _RAND_426 = {1{`RANDOM}};
  btb_426 = _RAND_426[31:0];
  _RAND_427 = {1{`RANDOM}};
  btb_427 = _RAND_427[31:0];
  _RAND_428 = {1{`RANDOM}};
  btb_428 = _RAND_428[31:0];
  _RAND_429 = {1{`RANDOM}};
  btb_429 = _RAND_429[31:0];
  _RAND_430 = {1{`RANDOM}};
  btb_430 = _RAND_430[31:0];
  _RAND_431 = {1{`RANDOM}};
  btb_431 = _RAND_431[31:0];
  _RAND_432 = {1{`RANDOM}};
  btb_432 = _RAND_432[31:0];
  _RAND_433 = {1{`RANDOM}};
  btb_433 = _RAND_433[31:0];
  _RAND_434 = {1{`RANDOM}};
  btb_434 = _RAND_434[31:0];
  _RAND_435 = {1{`RANDOM}};
  btb_435 = _RAND_435[31:0];
  _RAND_436 = {1{`RANDOM}};
  btb_436 = _RAND_436[31:0];
  _RAND_437 = {1{`RANDOM}};
  btb_437 = _RAND_437[31:0];
  _RAND_438 = {1{`RANDOM}};
  btb_438 = _RAND_438[31:0];
  _RAND_439 = {1{`RANDOM}};
  btb_439 = _RAND_439[31:0];
  _RAND_440 = {1{`RANDOM}};
  btb_440 = _RAND_440[31:0];
  _RAND_441 = {1{`RANDOM}};
  btb_441 = _RAND_441[31:0];
  _RAND_442 = {1{`RANDOM}};
  btb_442 = _RAND_442[31:0];
  _RAND_443 = {1{`RANDOM}};
  btb_443 = _RAND_443[31:0];
  _RAND_444 = {1{`RANDOM}};
  btb_444 = _RAND_444[31:0];
  _RAND_445 = {1{`RANDOM}};
  btb_445 = _RAND_445[31:0];
  _RAND_446 = {1{`RANDOM}};
  btb_446 = _RAND_446[31:0];
  _RAND_447 = {1{`RANDOM}};
  btb_447 = _RAND_447[31:0];
  _RAND_448 = {1{`RANDOM}};
  btb_448 = _RAND_448[31:0];
  _RAND_449 = {1{`RANDOM}};
  btb_449 = _RAND_449[31:0];
  _RAND_450 = {1{`RANDOM}};
  btb_450 = _RAND_450[31:0];
  _RAND_451 = {1{`RANDOM}};
  btb_451 = _RAND_451[31:0];
  _RAND_452 = {1{`RANDOM}};
  btb_452 = _RAND_452[31:0];
  _RAND_453 = {1{`RANDOM}};
  btb_453 = _RAND_453[31:0];
  _RAND_454 = {1{`RANDOM}};
  btb_454 = _RAND_454[31:0];
  _RAND_455 = {1{`RANDOM}};
  btb_455 = _RAND_455[31:0];
  _RAND_456 = {1{`RANDOM}};
  btb_456 = _RAND_456[31:0];
  _RAND_457 = {1{`RANDOM}};
  btb_457 = _RAND_457[31:0];
  _RAND_458 = {1{`RANDOM}};
  btb_458 = _RAND_458[31:0];
  _RAND_459 = {1{`RANDOM}};
  btb_459 = _RAND_459[31:0];
  _RAND_460 = {1{`RANDOM}};
  btb_460 = _RAND_460[31:0];
  _RAND_461 = {1{`RANDOM}};
  btb_461 = _RAND_461[31:0];
  _RAND_462 = {1{`RANDOM}};
  btb_462 = _RAND_462[31:0];
  _RAND_463 = {1{`RANDOM}};
  btb_463 = _RAND_463[31:0];
  _RAND_464 = {1{`RANDOM}};
  btb_464 = _RAND_464[31:0];
  _RAND_465 = {1{`RANDOM}};
  btb_465 = _RAND_465[31:0];
  _RAND_466 = {1{`RANDOM}};
  btb_466 = _RAND_466[31:0];
  _RAND_467 = {1{`RANDOM}};
  btb_467 = _RAND_467[31:0];
  _RAND_468 = {1{`RANDOM}};
  btb_468 = _RAND_468[31:0];
  _RAND_469 = {1{`RANDOM}};
  btb_469 = _RAND_469[31:0];
  _RAND_470 = {1{`RANDOM}};
  btb_470 = _RAND_470[31:0];
  _RAND_471 = {1{`RANDOM}};
  btb_471 = _RAND_471[31:0];
  _RAND_472 = {1{`RANDOM}};
  btb_472 = _RAND_472[31:0];
  _RAND_473 = {1{`RANDOM}};
  btb_473 = _RAND_473[31:0];
  _RAND_474 = {1{`RANDOM}};
  btb_474 = _RAND_474[31:0];
  _RAND_475 = {1{`RANDOM}};
  btb_475 = _RAND_475[31:0];
  _RAND_476 = {1{`RANDOM}};
  btb_476 = _RAND_476[31:0];
  _RAND_477 = {1{`RANDOM}};
  btb_477 = _RAND_477[31:0];
  _RAND_478 = {1{`RANDOM}};
  btb_478 = _RAND_478[31:0];
  _RAND_479 = {1{`RANDOM}};
  btb_479 = _RAND_479[31:0];
  _RAND_480 = {1{`RANDOM}};
  btb_480 = _RAND_480[31:0];
  _RAND_481 = {1{`RANDOM}};
  btb_481 = _RAND_481[31:0];
  _RAND_482 = {1{`RANDOM}};
  btb_482 = _RAND_482[31:0];
  _RAND_483 = {1{`RANDOM}};
  btb_483 = _RAND_483[31:0];
  _RAND_484 = {1{`RANDOM}};
  btb_484 = _RAND_484[31:0];
  _RAND_485 = {1{`RANDOM}};
  btb_485 = _RAND_485[31:0];
  _RAND_486 = {1{`RANDOM}};
  btb_486 = _RAND_486[31:0];
  _RAND_487 = {1{`RANDOM}};
  btb_487 = _RAND_487[31:0];
  _RAND_488 = {1{`RANDOM}};
  btb_488 = _RAND_488[31:0];
  _RAND_489 = {1{`RANDOM}};
  btb_489 = _RAND_489[31:0];
  _RAND_490 = {1{`RANDOM}};
  btb_490 = _RAND_490[31:0];
  _RAND_491 = {1{`RANDOM}};
  btb_491 = _RAND_491[31:0];
  _RAND_492 = {1{`RANDOM}};
  btb_492 = _RAND_492[31:0];
  _RAND_493 = {1{`RANDOM}};
  btb_493 = _RAND_493[31:0];
  _RAND_494 = {1{`RANDOM}};
  btb_494 = _RAND_494[31:0];
  _RAND_495 = {1{`RANDOM}};
  btb_495 = _RAND_495[31:0];
  _RAND_496 = {1{`RANDOM}};
  btb_496 = _RAND_496[31:0];
  _RAND_497 = {1{`RANDOM}};
  btb_497 = _RAND_497[31:0];
  _RAND_498 = {1{`RANDOM}};
  btb_498 = _RAND_498[31:0];
  _RAND_499 = {1{`RANDOM}};
  btb_499 = _RAND_499[31:0];
  _RAND_500 = {1{`RANDOM}};
  btb_500 = _RAND_500[31:0];
  _RAND_501 = {1{`RANDOM}};
  btb_501 = _RAND_501[31:0];
  _RAND_502 = {1{`RANDOM}};
  btb_502 = _RAND_502[31:0];
  _RAND_503 = {1{`RANDOM}};
  btb_503 = _RAND_503[31:0];
  _RAND_504 = {1{`RANDOM}};
  btb_504 = _RAND_504[31:0];
  _RAND_505 = {1{`RANDOM}};
  btb_505 = _RAND_505[31:0];
  _RAND_506 = {1{`RANDOM}};
  btb_506 = _RAND_506[31:0];
  _RAND_507 = {1{`RANDOM}};
  btb_507 = _RAND_507[31:0];
  _RAND_508 = {1{`RANDOM}};
  btb_508 = _RAND_508[31:0];
  _RAND_509 = {1{`RANDOM}};
  btb_509 = _RAND_509[31:0];
  _RAND_510 = {1{`RANDOM}};
  btb_510 = _RAND_510[31:0];
  _RAND_511 = {1{`RANDOM}};
  btb_511 = _RAND_511[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    btb_0 = 32'h0;
  end
  if (reset) begin
    btb_1 = 32'h0;
  end
  if (reset) begin
    btb_2 = 32'h0;
  end
  if (reset) begin
    btb_3 = 32'h0;
  end
  if (reset) begin
    btb_4 = 32'h0;
  end
  if (reset) begin
    btb_5 = 32'h0;
  end
  if (reset) begin
    btb_6 = 32'h0;
  end
  if (reset) begin
    btb_7 = 32'h0;
  end
  if (reset) begin
    btb_8 = 32'h0;
  end
  if (reset) begin
    btb_9 = 32'h0;
  end
  if (reset) begin
    btb_10 = 32'h0;
  end
  if (reset) begin
    btb_11 = 32'h0;
  end
  if (reset) begin
    btb_12 = 32'h0;
  end
  if (reset) begin
    btb_13 = 32'h0;
  end
  if (reset) begin
    btb_14 = 32'h0;
  end
  if (reset) begin
    btb_15 = 32'h0;
  end
  if (reset) begin
    btb_16 = 32'h0;
  end
  if (reset) begin
    btb_17 = 32'h0;
  end
  if (reset) begin
    btb_18 = 32'h0;
  end
  if (reset) begin
    btb_19 = 32'h0;
  end
  if (reset) begin
    btb_20 = 32'h0;
  end
  if (reset) begin
    btb_21 = 32'h0;
  end
  if (reset) begin
    btb_22 = 32'h0;
  end
  if (reset) begin
    btb_23 = 32'h0;
  end
  if (reset) begin
    btb_24 = 32'h0;
  end
  if (reset) begin
    btb_25 = 32'h0;
  end
  if (reset) begin
    btb_26 = 32'h0;
  end
  if (reset) begin
    btb_27 = 32'h0;
  end
  if (reset) begin
    btb_28 = 32'h0;
  end
  if (reset) begin
    btb_29 = 32'h0;
  end
  if (reset) begin
    btb_30 = 32'h0;
  end
  if (reset) begin
    btb_31 = 32'h0;
  end
  if (reset) begin
    btb_32 = 32'h0;
  end
  if (reset) begin
    btb_33 = 32'h0;
  end
  if (reset) begin
    btb_34 = 32'h0;
  end
  if (reset) begin
    btb_35 = 32'h0;
  end
  if (reset) begin
    btb_36 = 32'h0;
  end
  if (reset) begin
    btb_37 = 32'h0;
  end
  if (reset) begin
    btb_38 = 32'h0;
  end
  if (reset) begin
    btb_39 = 32'h0;
  end
  if (reset) begin
    btb_40 = 32'h0;
  end
  if (reset) begin
    btb_41 = 32'h0;
  end
  if (reset) begin
    btb_42 = 32'h0;
  end
  if (reset) begin
    btb_43 = 32'h0;
  end
  if (reset) begin
    btb_44 = 32'h0;
  end
  if (reset) begin
    btb_45 = 32'h0;
  end
  if (reset) begin
    btb_46 = 32'h0;
  end
  if (reset) begin
    btb_47 = 32'h0;
  end
  if (reset) begin
    btb_48 = 32'h0;
  end
  if (reset) begin
    btb_49 = 32'h0;
  end
  if (reset) begin
    btb_50 = 32'h0;
  end
  if (reset) begin
    btb_51 = 32'h0;
  end
  if (reset) begin
    btb_52 = 32'h0;
  end
  if (reset) begin
    btb_53 = 32'h0;
  end
  if (reset) begin
    btb_54 = 32'h0;
  end
  if (reset) begin
    btb_55 = 32'h0;
  end
  if (reset) begin
    btb_56 = 32'h0;
  end
  if (reset) begin
    btb_57 = 32'h0;
  end
  if (reset) begin
    btb_58 = 32'h0;
  end
  if (reset) begin
    btb_59 = 32'h0;
  end
  if (reset) begin
    btb_60 = 32'h0;
  end
  if (reset) begin
    btb_61 = 32'h0;
  end
  if (reset) begin
    btb_62 = 32'h0;
  end
  if (reset) begin
    btb_63 = 32'h0;
  end
  if (reset) begin
    btb_64 = 32'h0;
  end
  if (reset) begin
    btb_65 = 32'h0;
  end
  if (reset) begin
    btb_66 = 32'h0;
  end
  if (reset) begin
    btb_67 = 32'h0;
  end
  if (reset) begin
    btb_68 = 32'h0;
  end
  if (reset) begin
    btb_69 = 32'h0;
  end
  if (reset) begin
    btb_70 = 32'h0;
  end
  if (reset) begin
    btb_71 = 32'h0;
  end
  if (reset) begin
    btb_72 = 32'h0;
  end
  if (reset) begin
    btb_73 = 32'h0;
  end
  if (reset) begin
    btb_74 = 32'h0;
  end
  if (reset) begin
    btb_75 = 32'h0;
  end
  if (reset) begin
    btb_76 = 32'h0;
  end
  if (reset) begin
    btb_77 = 32'h0;
  end
  if (reset) begin
    btb_78 = 32'h0;
  end
  if (reset) begin
    btb_79 = 32'h0;
  end
  if (reset) begin
    btb_80 = 32'h0;
  end
  if (reset) begin
    btb_81 = 32'h0;
  end
  if (reset) begin
    btb_82 = 32'h0;
  end
  if (reset) begin
    btb_83 = 32'h0;
  end
  if (reset) begin
    btb_84 = 32'h0;
  end
  if (reset) begin
    btb_85 = 32'h0;
  end
  if (reset) begin
    btb_86 = 32'h0;
  end
  if (reset) begin
    btb_87 = 32'h0;
  end
  if (reset) begin
    btb_88 = 32'h0;
  end
  if (reset) begin
    btb_89 = 32'h0;
  end
  if (reset) begin
    btb_90 = 32'h0;
  end
  if (reset) begin
    btb_91 = 32'h0;
  end
  if (reset) begin
    btb_92 = 32'h0;
  end
  if (reset) begin
    btb_93 = 32'h0;
  end
  if (reset) begin
    btb_94 = 32'h0;
  end
  if (reset) begin
    btb_95 = 32'h0;
  end
  if (reset) begin
    btb_96 = 32'h0;
  end
  if (reset) begin
    btb_97 = 32'h0;
  end
  if (reset) begin
    btb_98 = 32'h0;
  end
  if (reset) begin
    btb_99 = 32'h0;
  end
  if (reset) begin
    btb_100 = 32'h0;
  end
  if (reset) begin
    btb_101 = 32'h0;
  end
  if (reset) begin
    btb_102 = 32'h0;
  end
  if (reset) begin
    btb_103 = 32'h0;
  end
  if (reset) begin
    btb_104 = 32'h0;
  end
  if (reset) begin
    btb_105 = 32'h0;
  end
  if (reset) begin
    btb_106 = 32'h0;
  end
  if (reset) begin
    btb_107 = 32'h0;
  end
  if (reset) begin
    btb_108 = 32'h0;
  end
  if (reset) begin
    btb_109 = 32'h0;
  end
  if (reset) begin
    btb_110 = 32'h0;
  end
  if (reset) begin
    btb_111 = 32'h0;
  end
  if (reset) begin
    btb_112 = 32'h0;
  end
  if (reset) begin
    btb_113 = 32'h0;
  end
  if (reset) begin
    btb_114 = 32'h0;
  end
  if (reset) begin
    btb_115 = 32'h0;
  end
  if (reset) begin
    btb_116 = 32'h0;
  end
  if (reset) begin
    btb_117 = 32'h0;
  end
  if (reset) begin
    btb_118 = 32'h0;
  end
  if (reset) begin
    btb_119 = 32'h0;
  end
  if (reset) begin
    btb_120 = 32'h0;
  end
  if (reset) begin
    btb_121 = 32'h0;
  end
  if (reset) begin
    btb_122 = 32'h0;
  end
  if (reset) begin
    btb_123 = 32'h0;
  end
  if (reset) begin
    btb_124 = 32'h0;
  end
  if (reset) begin
    btb_125 = 32'h0;
  end
  if (reset) begin
    btb_126 = 32'h0;
  end
  if (reset) begin
    btb_127 = 32'h0;
  end
  if (reset) begin
    btb_128 = 32'h0;
  end
  if (reset) begin
    btb_129 = 32'h0;
  end
  if (reset) begin
    btb_130 = 32'h0;
  end
  if (reset) begin
    btb_131 = 32'h0;
  end
  if (reset) begin
    btb_132 = 32'h0;
  end
  if (reset) begin
    btb_133 = 32'h0;
  end
  if (reset) begin
    btb_134 = 32'h0;
  end
  if (reset) begin
    btb_135 = 32'h0;
  end
  if (reset) begin
    btb_136 = 32'h0;
  end
  if (reset) begin
    btb_137 = 32'h0;
  end
  if (reset) begin
    btb_138 = 32'h0;
  end
  if (reset) begin
    btb_139 = 32'h0;
  end
  if (reset) begin
    btb_140 = 32'h0;
  end
  if (reset) begin
    btb_141 = 32'h0;
  end
  if (reset) begin
    btb_142 = 32'h0;
  end
  if (reset) begin
    btb_143 = 32'h0;
  end
  if (reset) begin
    btb_144 = 32'h0;
  end
  if (reset) begin
    btb_145 = 32'h0;
  end
  if (reset) begin
    btb_146 = 32'h0;
  end
  if (reset) begin
    btb_147 = 32'h0;
  end
  if (reset) begin
    btb_148 = 32'h0;
  end
  if (reset) begin
    btb_149 = 32'h0;
  end
  if (reset) begin
    btb_150 = 32'h0;
  end
  if (reset) begin
    btb_151 = 32'h0;
  end
  if (reset) begin
    btb_152 = 32'h0;
  end
  if (reset) begin
    btb_153 = 32'h0;
  end
  if (reset) begin
    btb_154 = 32'h0;
  end
  if (reset) begin
    btb_155 = 32'h0;
  end
  if (reset) begin
    btb_156 = 32'h0;
  end
  if (reset) begin
    btb_157 = 32'h0;
  end
  if (reset) begin
    btb_158 = 32'h0;
  end
  if (reset) begin
    btb_159 = 32'h0;
  end
  if (reset) begin
    btb_160 = 32'h0;
  end
  if (reset) begin
    btb_161 = 32'h0;
  end
  if (reset) begin
    btb_162 = 32'h0;
  end
  if (reset) begin
    btb_163 = 32'h0;
  end
  if (reset) begin
    btb_164 = 32'h0;
  end
  if (reset) begin
    btb_165 = 32'h0;
  end
  if (reset) begin
    btb_166 = 32'h0;
  end
  if (reset) begin
    btb_167 = 32'h0;
  end
  if (reset) begin
    btb_168 = 32'h0;
  end
  if (reset) begin
    btb_169 = 32'h0;
  end
  if (reset) begin
    btb_170 = 32'h0;
  end
  if (reset) begin
    btb_171 = 32'h0;
  end
  if (reset) begin
    btb_172 = 32'h0;
  end
  if (reset) begin
    btb_173 = 32'h0;
  end
  if (reset) begin
    btb_174 = 32'h0;
  end
  if (reset) begin
    btb_175 = 32'h0;
  end
  if (reset) begin
    btb_176 = 32'h0;
  end
  if (reset) begin
    btb_177 = 32'h0;
  end
  if (reset) begin
    btb_178 = 32'h0;
  end
  if (reset) begin
    btb_179 = 32'h0;
  end
  if (reset) begin
    btb_180 = 32'h0;
  end
  if (reset) begin
    btb_181 = 32'h0;
  end
  if (reset) begin
    btb_182 = 32'h0;
  end
  if (reset) begin
    btb_183 = 32'h0;
  end
  if (reset) begin
    btb_184 = 32'h0;
  end
  if (reset) begin
    btb_185 = 32'h0;
  end
  if (reset) begin
    btb_186 = 32'h0;
  end
  if (reset) begin
    btb_187 = 32'h0;
  end
  if (reset) begin
    btb_188 = 32'h0;
  end
  if (reset) begin
    btb_189 = 32'h0;
  end
  if (reset) begin
    btb_190 = 32'h0;
  end
  if (reset) begin
    btb_191 = 32'h0;
  end
  if (reset) begin
    btb_192 = 32'h0;
  end
  if (reset) begin
    btb_193 = 32'h0;
  end
  if (reset) begin
    btb_194 = 32'h0;
  end
  if (reset) begin
    btb_195 = 32'h0;
  end
  if (reset) begin
    btb_196 = 32'h0;
  end
  if (reset) begin
    btb_197 = 32'h0;
  end
  if (reset) begin
    btb_198 = 32'h0;
  end
  if (reset) begin
    btb_199 = 32'h0;
  end
  if (reset) begin
    btb_200 = 32'h0;
  end
  if (reset) begin
    btb_201 = 32'h0;
  end
  if (reset) begin
    btb_202 = 32'h0;
  end
  if (reset) begin
    btb_203 = 32'h0;
  end
  if (reset) begin
    btb_204 = 32'h0;
  end
  if (reset) begin
    btb_205 = 32'h0;
  end
  if (reset) begin
    btb_206 = 32'h0;
  end
  if (reset) begin
    btb_207 = 32'h0;
  end
  if (reset) begin
    btb_208 = 32'h0;
  end
  if (reset) begin
    btb_209 = 32'h0;
  end
  if (reset) begin
    btb_210 = 32'h0;
  end
  if (reset) begin
    btb_211 = 32'h0;
  end
  if (reset) begin
    btb_212 = 32'h0;
  end
  if (reset) begin
    btb_213 = 32'h0;
  end
  if (reset) begin
    btb_214 = 32'h0;
  end
  if (reset) begin
    btb_215 = 32'h0;
  end
  if (reset) begin
    btb_216 = 32'h0;
  end
  if (reset) begin
    btb_217 = 32'h0;
  end
  if (reset) begin
    btb_218 = 32'h0;
  end
  if (reset) begin
    btb_219 = 32'h0;
  end
  if (reset) begin
    btb_220 = 32'h0;
  end
  if (reset) begin
    btb_221 = 32'h0;
  end
  if (reset) begin
    btb_222 = 32'h0;
  end
  if (reset) begin
    btb_223 = 32'h0;
  end
  if (reset) begin
    btb_224 = 32'h0;
  end
  if (reset) begin
    btb_225 = 32'h0;
  end
  if (reset) begin
    btb_226 = 32'h0;
  end
  if (reset) begin
    btb_227 = 32'h0;
  end
  if (reset) begin
    btb_228 = 32'h0;
  end
  if (reset) begin
    btb_229 = 32'h0;
  end
  if (reset) begin
    btb_230 = 32'h0;
  end
  if (reset) begin
    btb_231 = 32'h0;
  end
  if (reset) begin
    btb_232 = 32'h0;
  end
  if (reset) begin
    btb_233 = 32'h0;
  end
  if (reset) begin
    btb_234 = 32'h0;
  end
  if (reset) begin
    btb_235 = 32'h0;
  end
  if (reset) begin
    btb_236 = 32'h0;
  end
  if (reset) begin
    btb_237 = 32'h0;
  end
  if (reset) begin
    btb_238 = 32'h0;
  end
  if (reset) begin
    btb_239 = 32'h0;
  end
  if (reset) begin
    btb_240 = 32'h0;
  end
  if (reset) begin
    btb_241 = 32'h0;
  end
  if (reset) begin
    btb_242 = 32'h0;
  end
  if (reset) begin
    btb_243 = 32'h0;
  end
  if (reset) begin
    btb_244 = 32'h0;
  end
  if (reset) begin
    btb_245 = 32'h0;
  end
  if (reset) begin
    btb_246 = 32'h0;
  end
  if (reset) begin
    btb_247 = 32'h0;
  end
  if (reset) begin
    btb_248 = 32'h0;
  end
  if (reset) begin
    btb_249 = 32'h0;
  end
  if (reset) begin
    btb_250 = 32'h0;
  end
  if (reset) begin
    btb_251 = 32'h0;
  end
  if (reset) begin
    btb_252 = 32'h0;
  end
  if (reset) begin
    btb_253 = 32'h0;
  end
  if (reset) begin
    btb_254 = 32'h0;
  end
  if (reset) begin
    btb_255 = 32'h0;
  end
  if (reset) begin
    btb_256 = 32'h0;
  end
  if (reset) begin
    btb_257 = 32'h0;
  end
  if (reset) begin
    btb_258 = 32'h0;
  end
  if (reset) begin
    btb_259 = 32'h0;
  end
  if (reset) begin
    btb_260 = 32'h0;
  end
  if (reset) begin
    btb_261 = 32'h0;
  end
  if (reset) begin
    btb_262 = 32'h0;
  end
  if (reset) begin
    btb_263 = 32'h0;
  end
  if (reset) begin
    btb_264 = 32'h0;
  end
  if (reset) begin
    btb_265 = 32'h0;
  end
  if (reset) begin
    btb_266 = 32'h0;
  end
  if (reset) begin
    btb_267 = 32'h0;
  end
  if (reset) begin
    btb_268 = 32'h0;
  end
  if (reset) begin
    btb_269 = 32'h0;
  end
  if (reset) begin
    btb_270 = 32'h0;
  end
  if (reset) begin
    btb_271 = 32'h0;
  end
  if (reset) begin
    btb_272 = 32'h0;
  end
  if (reset) begin
    btb_273 = 32'h0;
  end
  if (reset) begin
    btb_274 = 32'h0;
  end
  if (reset) begin
    btb_275 = 32'h0;
  end
  if (reset) begin
    btb_276 = 32'h0;
  end
  if (reset) begin
    btb_277 = 32'h0;
  end
  if (reset) begin
    btb_278 = 32'h0;
  end
  if (reset) begin
    btb_279 = 32'h0;
  end
  if (reset) begin
    btb_280 = 32'h0;
  end
  if (reset) begin
    btb_281 = 32'h0;
  end
  if (reset) begin
    btb_282 = 32'h0;
  end
  if (reset) begin
    btb_283 = 32'h0;
  end
  if (reset) begin
    btb_284 = 32'h0;
  end
  if (reset) begin
    btb_285 = 32'h0;
  end
  if (reset) begin
    btb_286 = 32'h0;
  end
  if (reset) begin
    btb_287 = 32'h0;
  end
  if (reset) begin
    btb_288 = 32'h0;
  end
  if (reset) begin
    btb_289 = 32'h0;
  end
  if (reset) begin
    btb_290 = 32'h0;
  end
  if (reset) begin
    btb_291 = 32'h0;
  end
  if (reset) begin
    btb_292 = 32'h0;
  end
  if (reset) begin
    btb_293 = 32'h0;
  end
  if (reset) begin
    btb_294 = 32'h0;
  end
  if (reset) begin
    btb_295 = 32'h0;
  end
  if (reset) begin
    btb_296 = 32'h0;
  end
  if (reset) begin
    btb_297 = 32'h0;
  end
  if (reset) begin
    btb_298 = 32'h0;
  end
  if (reset) begin
    btb_299 = 32'h0;
  end
  if (reset) begin
    btb_300 = 32'h0;
  end
  if (reset) begin
    btb_301 = 32'h0;
  end
  if (reset) begin
    btb_302 = 32'h0;
  end
  if (reset) begin
    btb_303 = 32'h0;
  end
  if (reset) begin
    btb_304 = 32'h0;
  end
  if (reset) begin
    btb_305 = 32'h0;
  end
  if (reset) begin
    btb_306 = 32'h0;
  end
  if (reset) begin
    btb_307 = 32'h0;
  end
  if (reset) begin
    btb_308 = 32'h0;
  end
  if (reset) begin
    btb_309 = 32'h0;
  end
  if (reset) begin
    btb_310 = 32'h0;
  end
  if (reset) begin
    btb_311 = 32'h0;
  end
  if (reset) begin
    btb_312 = 32'h0;
  end
  if (reset) begin
    btb_313 = 32'h0;
  end
  if (reset) begin
    btb_314 = 32'h0;
  end
  if (reset) begin
    btb_315 = 32'h0;
  end
  if (reset) begin
    btb_316 = 32'h0;
  end
  if (reset) begin
    btb_317 = 32'h0;
  end
  if (reset) begin
    btb_318 = 32'h0;
  end
  if (reset) begin
    btb_319 = 32'h0;
  end
  if (reset) begin
    btb_320 = 32'h0;
  end
  if (reset) begin
    btb_321 = 32'h0;
  end
  if (reset) begin
    btb_322 = 32'h0;
  end
  if (reset) begin
    btb_323 = 32'h0;
  end
  if (reset) begin
    btb_324 = 32'h0;
  end
  if (reset) begin
    btb_325 = 32'h0;
  end
  if (reset) begin
    btb_326 = 32'h0;
  end
  if (reset) begin
    btb_327 = 32'h0;
  end
  if (reset) begin
    btb_328 = 32'h0;
  end
  if (reset) begin
    btb_329 = 32'h0;
  end
  if (reset) begin
    btb_330 = 32'h0;
  end
  if (reset) begin
    btb_331 = 32'h0;
  end
  if (reset) begin
    btb_332 = 32'h0;
  end
  if (reset) begin
    btb_333 = 32'h0;
  end
  if (reset) begin
    btb_334 = 32'h0;
  end
  if (reset) begin
    btb_335 = 32'h0;
  end
  if (reset) begin
    btb_336 = 32'h0;
  end
  if (reset) begin
    btb_337 = 32'h0;
  end
  if (reset) begin
    btb_338 = 32'h0;
  end
  if (reset) begin
    btb_339 = 32'h0;
  end
  if (reset) begin
    btb_340 = 32'h0;
  end
  if (reset) begin
    btb_341 = 32'h0;
  end
  if (reset) begin
    btb_342 = 32'h0;
  end
  if (reset) begin
    btb_343 = 32'h0;
  end
  if (reset) begin
    btb_344 = 32'h0;
  end
  if (reset) begin
    btb_345 = 32'h0;
  end
  if (reset) begin
    btb_346 = 32'h0;
  end
  if (reset) begin
    btb_347 = 32'h0;
  end
  if (reset) begin
    btb_348 = 32'h0;
  end
  if (reset) begin
    btb_349 = 32'h0;
  end
  if (reset) begin
    btb_350 = 32'h0;
  end
  if (reset) begin
    btb_351 = 32'h0;
  end
  if (reset) begin
    btb_352 = 32'h0;
  end
  if (reset) begin
    btb_353 = 32'h0;
  end
  if (reset) begin
    btb_354 = 32'h0;
  end
  if (reset) begin
    btb_355 = 32'h0;
  end
  if (reset) begin
    btb_356 = 32'h0;
  end
  if (reset) begin
    btb_357 = 32'h0;
  end
  if (reset) begin
    btb_358 = 32'h0;
  end
  if (reset) begin
    btb_359 = 32'h0;
  end
  if (reset) begin
    btb_360 = 32'h0;
  end
  if (reset) begin
    btb_361 = 32'h0;
  end
  if (reset) begin
    btb_362 = 32'h0;
  end
  if (reset) begin
    btb_363 = 32'h0;
  end
  if (reset) begin
    btb_364 = 32'h0;
  end
  if (reset) begin
    btb_365 = 32'h0;
  end
  if (reset) begin
    btb_366 = 32'h0;
  end
  if (reset) begin
    btb_367 = 32'h0;
  end
  if (reset) begin
    btb_368 = 32'h0;
  end
  if (reset) begin
    btb_369 = 32'h0;
  end
  if (reset) begin
    btb_370 = 32'h0;
  end
  if (reset) begin
    btb_371 = 32'h0;
  end
  if (reset) begin
    btb_372 = 32'h0;
  end
  if (reset) begin
    btb_373 = 32'h0;
  end
  if (reset) begin
    btb_374 = 32'h0;
  end
  if (reset) begin
    btb_375 = 32'h0;
  end
  if (reset) begin
    btb_376 = 32'h0;
  end
  if (reset) begin
    btb_377 = 32'h0;
  end
  if (reset) begin
    btb_378 = 32'h0;
  end
  if (reset) begin
    btb_379 = 32'h0;
  end
  if (reset) begin
    btb_380 = 32'h0;
  end
  if (reset) begin
    btb_381 = 32'h0;
  end
  if (reset) begin
    btb_382 = 32'h0;
  end
  if (reset) begin
    btb_383 = 32'h0;
  end
  if (reset) begin
    btb_384 = 32'h0;
  end
  if (reset) begin
    btb_385 = 32'h0;
  end
  if (reset) begin
    btb_386 = 32'h0;
  end
  if (reset) begin
    btb_387 = 32'h0;
  end
  if (reset) begin
    btb_388 = 32'h0;
  end
  if (reset) begin
    btb_389 = 32'h0;
  end
  if (reset) begin
    btb_390 = 32'h0;
  end
  if (reset) begin
    btb_391 = 32'h0;
  end
  if (reset) begin
    btb_392 = 32'h0;
  end
  if (reset) begin
    btb_393 = 32'h0;
  end
  if (reset) begin
    btb_394 = 32'h0;
  end
  if (reset) begin
    btb_395 = 32'h0;
  end
  if (reset) begin
    btb_396 = 32'h0;
  end
  if (reset) begin
    btb_397 = 32'h0;
  end
  if (reset) begin
    btb_398 = 32'h0;
  end
  if (reset) begin
    btb_399 = 32'h0;
  end
  if (reset) begin
    btb_400 = 32'h0;
  end
  if (reset) begin
    btb_401 = 32'h0;
  end
  if (reset) begin
    btb_402 = 32'h0;
  end
  if (reset) begin
    btb_403 = 32'h0;
  end
  if (reset) begin
    btb_404 = 32'h0;
  end
  if (reset) begin
    btb_405 = 32'h0;
  end
  if (reset) begin
    btb_406 = 32'h0;
  end
  if (reset) begin
    btb_407 = 32'h0;
  end
  if (reset) begin
    btb_408 = 32'h0;
  end
  if (reset) begin
    btb_409 = 32'h0;
  end
  if (reset) begin
    btb_410 = 32'h0;
  end
  if (reset) begin
    btb_411 = 32'h0;
  end
  if (reset) begin
    btb_412 = 32'h0;
  end
  if (reset) begin
    btb_413 = 32'h0;
  end
  if (reset) begin
    btb_414 = 32'h0;
  end
  if (reset) begin
    btb_415 = 32'h0;
  end
  if (reset) begin
    btb_416 = 32'h0;
  end
  if (reset) begin
    btb_417 = 32'h0;
  end
  if (reset) begin
    btb_418 = 32'h0;
  end
  if (reset) begin
    btb_419 = 32'h0;
  end
  if (reset) begin
    btb_420 = 32'h0;
  end
  if (reset) begin
    btb_421 = 32'h0;
  end
  if (reset) begin
    btb_422 = 32'h0;
  end
  if (reset) begin
    btb_423 = 32'h0;
  end
  if (reset) begin
    btb_424 = 32'h0;
  end
  if (reset) begin
    btb_425 = 32'h0;
  end
  if (reset) begin
    btb_426 = 32'h0;
  end
  if (reset) begin
    btb_427 = 32'h0;
  end
  if (reset) begin
    btb_428 = 32'h0;
  end
  if (reset) begin
    btb_429 = 32'h0;
  end
  if (reset) begin
    btb_430 = 32'h0;
  end
  if (reset) begin
    btb_431 = 32'h0;
  end
  if (reset) begin
    btb_432 = 32'h0;
  end
  if (reset) begin
    btb_433 = 32'h0;
  end
  if (reset) begin
    btb_434 = 32'h0;
  end
  if (reset) begin
    btb_435 = 32'h0;
  end
  if (reset) begin
    btb_436 = 32'h0;
  end
  if (reset) begin
    btb_437 = 32'h0;
  end
  if (reset) begin
    btb_438 = 32'h0;
  end
  if (reset) begin
    btb_439 = 32'h0;
  end
  if (reset) begin
    btb_440 = 32'h0;
  end
  if (reset) begin
    btb_441 = 32'h0;
  end
  if (reset) begin
    btb_442 = 32'h0;
  end
  if (reset) begin
    btb_443 = 32'h0;
  end
  if (reset) begin
    btb_444 = 32'h0;
  end
  if (reset) begin
    btb_445 = 32'h0;
  end
  if (reset) begin
    btb_446 = 32'h0;
  end
  if (reset) begin
    btb_447 = 32'h0;
  end
  if (reset) begin
    btb_448 = 32'h0;
  end
  if (reset) begin
    btb_449 = 32'h0;
  end
  if (reset) begin
    btb_450 = 32'h0;
  end
  if (reset) begin
    btb_451 = 32'h0;
  end
  if (reset) begin
    btb_452 = 32'h0;
  end
  if (reset) begin
    btb_453 = 32'h0;
  end
  if (reset) begin
    btb_454 = 32'h0;
  end
  if (reset) begin
    btb_455 = 32'h0;
  end
  if (reset) begin
    btb_456 = 32'h0;
  end
  if (reset) begin
    btb_457 = 32'h0;
  end
  if (reset) begin
    btb_458 = 32'h0;
  end
  if (reset) begin
    btb_459 = 32'h0;
  end
  if (reset) begin
    btb_460 = 32'h0;
  end
  if (reset) begin
    btb_461 = 32'h0;
  end
  if (reset) begin
    btb_462 = 32'h0;
  end
  if (reset) begin
    btb_463 = 32'h0;
  end
  if (reset) begin
    btb_464 = 32'h0;
  end
  if (reset) begin
    btb_465 = 32'h0;
  end
  if (reset) begin
    btb_466 = 32'h0;
  end
  if (reset) begin
    btb_467 = 32'h0;
  end
  if (reset) begin
    btb_468 = 32'h0;
  end
  if (reset) begin
    btb_469 = 32'h0;
  end
  if (reset) begin
    btb_470 = 32'h0;
  end
  if (reset) begin
    btb_471 = 32'h0;
  end
  if (reset) begin
    btb_472 = 32'h0;
  end
  if (reset) begin
    btb_473 = 32'h0;
  end
  if (reset) begin
    btb_474 = 32'h0;
  end
  if (reset) begin
    btb_475 = 32'h0;
  end
  if (reset) begin
    btb_476 = 32'h0;
  end
  if (reset) begin
    btb_477 = 32'h0;
  end
  if (reset) begin
    btb_478 = 32'h0;
  end
  if (reset) begin
    btb_479 = 32'h0;
  end
  if (reset) begin
    btb_480 = 32'h0;
  end
  if (reset) begin
    btb_481 = 32'h0;
  end
  if (reset) begin
    btb_482 = 32'h0;
  end
  if (reset) begin
    btb_483 = 32'h0;
  end
  if (reset) begin
    btb_484 = 32'h0;
  end
  if (reset) begin
    btb_485 = 32'h0;
  end
  if (reset) begin
    btb_486 = 32'h0;
  end
  if (reset) begin
    btb_487 = 32'h0;
  end
  if (reset) begin
    btb_488 = 32'h0;
  end
  if (reset) begin
    btb_489 = 32'h0;
  end
  if (reset) begin
    btb_490 = 32'h0;
  end
  if (reset) begin
    btb_491 = 32'h0;
  end
  if (reset) begin
    btb_492 = 32'h0;
  end
  if (reset) begin
    btb_493 = 32'h0;
  end
  if (reset) begin
    btb_494 = 32'h0;
  end
  if (reset) begin
    btb_495 = 32'h0;
  end
  if (reset) begin
    btb_496 = 32'h0;
  end
  if (reset) begin
    btb_497 = 32'h0;
  end
  if (reset) begin
    btb_498 = 32'h0;
  end
  if (reset) begin
    btb_499 = 32'h0;
  end
  if (reset) begin
    btb_500 = 32'h0;
  end
  if (reset) begin
    btb_501 = 32'h0;
  end
  if (reset) begin
    btb_502 = 32'h0;
  end
  if (reset) begin
    btb_503 = 32'h0;
  end
  if (reset) begin
    btb_504 = 32'h0;
  end
  if (reset) begin
    btb_505 = 32'h0;
  end
  if (reset) begin
    btb_506 = 32'h0;
  end
  if (reset) begin
    btb_507 = 32'h0;
  end
  if (reset) begin
    btb_508 = 32'h0;
  end
  if (reset) begin
    btb_509 = 32'h0;
  end
  if (reset) begin
    btb_510 = 32'h0;
  end
  if (reset) begin
    btb_511 = 32'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module data_ram_simple_two_ports_36(
  input         clock,
  input         reset,
  input         io_wea,
  input  [8:0]  io_addra,
  input  [31:0] io_dina,
  input  [8:0]  io_addrb,
  output [31:0] io_doutb
);
  wire  Look_up_table_read_first__clock; // @[ip_user.scala 97:23]
  wire  Look_up_table_read_first__reset; // @[ip_user.scala 97:23]
  wire [8:0] Look_up_table_read_first__io_ar_addr; // @[ip_user.scala 97:23]
  wire [8:0] Look_up_table_read_first__io_aw_addr; // @[ip_user.scala 97:23]
  wire  Look_up_table_read_first__io_write; // @[ip_user.scala 97:23]
  wire [31:0] Look_up_table_read_first__io_in; // @[ip_user.scala 97:23]
  wire [31:0] Look_up_table_read_first__io_out; // @[ip_user.scala 97:23]
  Look_up_table_read_first__36 Look_up_table_read_first_ ( // @[ip_user.scala 97:23]
    .clock(Look_up_table_read_first__clock),
    .reset(Look_up_table_read_first__reset),
    .io_ar_addr(Look_up_table_read_first__io_ar_addr),
    .io_aw_addr(Look_up_table_read_first__io_aw_addr),
    .io_write(Look_up_table_read_first__io_write),
    .io_in(Look_up_table_read_first__io_in),
    .io_out(Look_up_table_read_first__io_out)
  );
  assign io_doutb = Look_up_table_read_first__io_out; // @[ip_user.scala 102:19]
  assign Look_up_table_read_first__clock = clock;
  assign Look_up_table_read_first__reset = reset;
  assign Look_up_table_read_first__io_ar_addr = io_addra; // @[ip_user.scala 98:19]
  assign Look_up_table_read_first__io_aw_addr = io_addrb; // @[ip_user.scala 99:19]
  assign Look_up_table_read_first__io_write = io_wea; // @[ip_user.scala 101:19]
  assign Look_up_table_read_first__io_in = io_dina; // @[ip_user.scala 100:19]
endmodule
module btb_data_with_block_ram(
  input         clock,
  input         reset,
  input         io_wen,
  input  [8:0]  io_raddr,
  input  [8:0]  io_waddr,
  input  [63:0] io_wdata,
  output [63:0] io_rdata
);
  wire  btb_data_ram_0_clock; // @[BTB.scala 189:32]
  wire  btb_data_ram_0_reset; // @[BTB.scala 189:32]
  wire  btb_data_ram_0_io_wea; // @[BTB.scala 189:32]
  wire [8:0] btb_data_ram_0_io_addra; // @[BTB.scala 189:32]
  wire [31:0] btb_data_ram_0_io_dina; // @[BTB.scala 189:32]
  wire [8:0] btb_data_ram_0_io_addrb; // @[BTB.scala 189:32]
  wire [31:0] btb_data_ram_0_io_doutb; // @[BTB.scala 189:32]
  data_ram_simple_two_ports_36 btb_data_ram_0 ( // @[BTB.scala 189:32]
    .clock(btb_data_ram_0_clock),
    .reset(btb_data_ram_0_reset),
    .io_wea(btb_data_ram_0_io_wea),
    .io_addra(btb_data_ram_0_io_addra),
    .io_dina(btb_data_ram_0_io_dina),
    .io_addrb(btb_data_ram_0_io_addrb),
    .io_doutb(btb_data_ram_0_io_doutb)
  );
  assign io_rdata = {{32'd0}, btb_data_ram_0_io_doutb}; // @[BTB.scala 198:18]
  assign btb_data_ram_0_clock = clock;
  assign btb_data_ram_0_reset = reset;
  assign btb_data_ram_0_io_wea = io_wen; // @[BTB.scala 194:28]
  assign btb_data_ram_0_io_addra = io_waddr; // @[BTB.scala 195:29]
  assign btb_data_ram_0_io_dina = io_wdata[31:0]; // @[BTB.scala 197:28]
  assign btb_data_ram_0_io_addrb = io_raddr; // @[BTB.scala 196:29]
endmodule
module BTB_banks_oneissue_with_block_ram(
  input         clock,
  input         reset,
  input  [63:0] io_ar_addr_L,
  input  [63:0] io_aw_addr,
  input  [63:0] io_aw_target_addr,
  input         io_write,
  output [63:0] io_out_L,
  output        io_hit_L
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  btb_tag_with_block_ram_clock; // @[BTB.scala 249:54]
  wire  btb_tag_with_block_ram_reset; // @[BTB.scala 249:54]
  wire  btb_tag_with_block_ram_io_wen; // @[BTB.scala 249:54]
  wire [8:0] btb_tag_with_block_ram_io_raddr; // @[BTB.scala 249:54]
  wire [8:0] btb_tag_with_block_ram_io_waddr; // @[BTB.scala 249:54]
  wire [7:0] btb_tag_with_block_ram_io_wdata; // @[BTB.scala 249:54]
  wire [7:0] btb_tag_with_block_ram_io_rdata; // @[BTB.scala 249:54]
  wire  btb_tag_with_block_ram_1_clock; // @[BTB.scala 249:54]
  wire  btb_tag_with_block_ram_1_reset; // @[BTB.scala 249:54]
  wire  btb_tag_with_block_ram_1_io_wen; // @[BTB.scala 249:54]
  wire [8:0] btb_tag_with_block_ram_1_io_raddr; // @[BTB.scala 249:54]
  wire [8:0] btb_tag_with_block_ram_1_io_waddr; // @[BTB.scala 249:54]
  wire [7:0] btb_tag_with_block_ram_1_io_wdata; // @[BTB.scala 249:54]
  wire [7:0] btb_tag_with_block_ram_1_io_rdata; // @[BTB.scala 249:54]
  wire  btb_tag_with_block_ram_2_clock; // @[BTB.scala 249:54]
  wire  btb_tag_with_block_ram_2_reset; // @[BTB.scala 249:54]
  wire  btb_tag_with_block_ram_2_io_wen; // @[BTB.scala 249:54]
  wire [8:0] btb_tag_with_block_ram_2_io_raddr; // @[BTB.scala 249:54]
  wire [8:0] btb_tag_with_block_ram_2_io_waddr; // @[BTB.scala 249:54]
  wire [7:0] btb_tag_with_block_ram_2_io_wdata; // @[BTB.scala 249:54]
  wire [7:0] btb_tag_with_block_ram_2_io_rdata; // @[BTB.scala 249:54]
  wire  btb_tag_with_block_ram_3_clock; // @[BTB.scala 249:54]
  wire  btb_tag_with_block_ram_3_reset; // @[BTB.scala 249:54]
  wire  btb_tag_with_block_ram_3_io_wen; // @[BTB.scala 249:54]
  wire [8:0] btb_tag_with_block_ram_3_io_raddr; // @[BTB.scala 249:54]
  wire [8:0] btb_tag_with_block_ram_3_io_waddr; // @[BTB.scala 249:54]
  wire [7:0] btb_tag_with_block_ram_3_io_wdata; // @[BTB.scala 249:54]
  wire [7:0] btb_tag_with_block_ram_3_io_rdata; // @[BTB.scala 249:54]
  wire  btb_data_with_block_ram_clock; // @[BTB.scala 250:54]
  wire  btb_data_with_block_ram_reset; // @[BTB.scala 250:54]
  wire  btb_data_with_block_ram_io_wen; // @[BTB.scala 250:54]
  wire [8:0] btb_data_with_block_ram_io_raddr; // @[BTB.scala 250:54]
  wire [8:0] btb_data_with_block_ram_io_waddr; // @[BTB.scala 250:54]
  wire [63:0] btb_data_with_block_ram_io_wdata; // @[BTB.scala 250:54]
  wire [63:0] btb_data_with_block_ram_io_rdata; // @[BTB.scala 250:54]
  wire  btb_data_with_block_ram_1_clock; // @[BTB.scala 250:54]
  wire  btb_data_with_block_ram_1_reset; // @[BTB.scala 250:54]
  wire  btb_data_with_block_ram_1_io_wen; // @[BTB.scala 250:54]
  wire [8:0] btb_data_with_block_ram_1_io_raddr; // @[BTB.scala 250:54]
  wire [8:0] btb_data_with_block_ram_1_io_waddr; // @[BTB.scala 250:54]
  wire [63:0] btb_data_with_block_ram_1_io_wdata; // @[BTB.scala 250:54]
  wire [63:0] btb_data_with_block_ram_1_io_rdata; // @[BTB.scala 250:54]
  wire  btb_data_with_block_ram_2_clock; // @[BTB.scala 250:54]
  wire  btb_data_with_block_ram_2_reset; // @[BTB.scala 250:54]
  wire  btb_data_with_block_ram_2_io_wen; // @[BTB.scala 250:54]
  wire [8:0] btb_data_with_block_ram_2_io_raddr; // @[BTB.scala 250:54]
  wire [8:0] btb_data_with_block_ram_2_io_waddr; // @[BTB.scala 250:54]
  wire [63:0] btb_data_with_block_ram_2_io_wdata; // @[BTB.scala 250:54]
  wire [63:0] btb_data_with_block_ram_2_io_rdata; // @[BTB.scala 250:54]
  wire  btb_data_with_block_ram_3_clock; // @[BTB.scala 250:54]
  wire  btb_data_with_block_ram_3_reset; // @[BTB.scala 250:54]
  wire  btb_data_with_block_ram_3_io_wen; // @[BTB.scala 250:54]
  wire [8:0] btb_data_with_block_ram_3_io_raddr; // @[BTB.scala 250:54]
  wire [8:0] btb_data_with_block_ram_3_io_waddr; // @[BTB.scala 250:54]
  wire [63:0] btb_data_with_block_ram_3_io_wdata; // @[BTB.scala 250:54]
  wire [63:0] btb_data_with_block_ram_3_io_rdata; // @[BTB.scala 250:54]
  wire  _btb_banks_0_wen_T_1 = io_aw_addr[3:2] == 2'h0; // @[BTB.scala 253:62]
  wire  _btb_banks_1_wen_T_1 = io_aw_addr[3:2] == 2'h1; // @[BTB.scala 253:62]
  wire  _btb_banks_2_wen_T_1 = io_aw_addr[3:2] == 2'h2; // @[BTB.scala 253:62]
  wire  _btb_banks_3_wen_T_1 = io_aw_addr[3:2] == 2'h3; // @[BTB.scala 253:62]
  reg [63:0] ar_addr_reg; // @[BTB.scala 263:30]
  wire [63:0] btb_banks_0_rdata = btb_data_with_block_ram_io_rdata; // @[BTB.scala 250:{28,28}]
  wire [63:0] btb_banks_1_rdata = btb_data_with_block_ram_1_io_rdata; // @[BTB.scala 250:{28,28}]
  wire [63:0] _GEN_1 = 2'h1 == ar_addr_reg[3:2] ? btb_banks_1_rdata : btb_banks_0_rdata; // @[BTB.scala 265:{14,14}]
  wire [63:0] btb_banks_2_rdata = btb_data_with_block_ram_2_io_rdata; // @[BTB.scala 250:{28,28}]
  wire [63:0] _GEN_2 = 2'h2 == ar_addr_reg[3:2] ? btb_banks_2_rdata : _GEN_1; // @[BTB.scala 265:{14,14}]
  wire [63:0] btb_banks_3_rdata = btb_data_with_block_ram_3_io_rdata; // @[BTB.scala 250:{28,28}]
  wire [4:0] _tag_banks_0_wdata_T_1 = {1'h1,io_aw_addr[16:13]}; // @[Cat.scala 31:58]
  wire [7:0] tag_banks_0_rdata = btb_tag_with_block_ram_io_rdata; // @[BTB.scala 249:{28,28}]
  wire [7:0] tag_banks_1_rdata = btb_tag_with_block_ram_1_io_rdata; // @[BTB.scala 249:{28,28}]
  wire [7:0] _GEN_13 = 2'h1 == ar_addr_reg[3:2] ? tag_banks_1_rdata : tag_banks_0_rdata; // @[BTB.scala 286:{67,67}]
  wire [7:0] tag_banks_2_rdata = btb_tag_with_block_ram_2_io_rdata; // @[BTB.scala 249:{28,28}]
  wire [7:0] _GEN_14 = 2'h2 == ar_addr_reg[3:2] ? tag_banks_2_rdata : _GEN_13; // @[BTB.scala 286:{67,67}]
  wire [7:0] tag_banks_3_rdata = btb_tag_with_block_ram_3_io_rdata; // @[BTB.scala 249:{28,28}]
  wire [7:0] _GEN_15 = 2'h3 == ar_addr_reg[3:2] ? tag_banks_3_rdata : _GEN_14; // @[BTB.scala 286:{67,67}]
  btb_tag_with_block_ram btb_tag_with_block_ram ( // @[BTB.scala 249:54]
    .clock(btb_tag_with_block_ram_clock),
    .reset(btb_tag_with_block_ram_reset),
    .io_wen(btb_tag_with_block_ram_io_wen),
    .io_raddr(btb_tag_with_block_ram_io_raddr),
    .io_waddr(btb_tag_with_block_ram_io_waddr),
    .io_wdata(btb_tag_with_block_ram_io_wdata),
    .io_rdata(btb_tag_with_block_ram_io_rdata)
  );
  btb_tag_with_block_ram btb_tag_with_block_ram_1 ( // @[BTB.scala 249:54]
    .clock(btb_tag_with_block_ram_1_clock),
    .reset(btb_tag_with_block_ram_1_reset),
    .io_wen(btb_tag_with_block_ram_1_io_wen),
    .io_raddr(btb_tag_with_block_ram_1_io_raddr),
    .io_waddr(btb_tag_with_block_ram_1_io_waddr),
    .io_wdata(btb_tag_with_block_ram_1_io_wdata),
    .io_rdata(btb_tag_with_block_ram_1_io_rdata)
  );
  btb_tag_with_block_ram btb_tag_with_block_ram_2 ( // @[BTB.scala 249:54]
    .clock(btb_tag_with_block_ram_2_clock),
    .reset(btb_tag_with_block_ram_2_reset),
    .io_wen(btb_tag_with_block_ram_2_io_wen),
    .io_raddr(btb_tag_with_block_ram_2_io_raddr),
    .io_waddr(btb_tag_with_block_ram_2_io_waddr),
    .io_wdata(btb_tag_with_block_ram_2_io_wdata),
    .io_rdata(btb_tag_with_block_ram_2_io_rdata)
  );
  btb_tag_with_block_ram btb_tag_with_block_ram_3 ( // @[BTB.scala 249:54]
    .clock(btb_tag_with_block_ram_3_clock),
    .reset(btb_tag_with_block_ram_3_reset),
    .io_wen(btb_tag_with_block_ram_3_io_wen),
    .io_raddr(btb_tag_with_block_ram_3_io_raddr),
    .io_waddr(btb_tag_with_block_ram_3_io_waddr),
    .io_wdata(btb_tag_with_block_ram_3_io_wdata),
    .io_rdata(btb_tag_with_block_ram_3_io_rdata)
  );
  btb_data_with_block_ram btb_data_with_block_ram ( // @[BTB.scala 250:54]
    .clock(btb_data_with_block_ram_clock),
    .reset(btb_data_with_block_ram_reset),
    .io_wen(btb_data_with_block_ram_io_wen),
    .io_raddr(btb_data_with_block_ram_io_raddr),
    .io_waddr(btb_data_with_block_ram_io_waddr),
    .io_wdata(btb_data_with_block_ram_io_wdata),
    .io_rdata(btb_data_with_block_ram_io_rdata)
  );
  btb_data_with_block_ram btb_data_with_block_ram_1 ( // @[BTB.scala 250:54]
    .clock(btb_data_with_block_ram_1_clock),
    .reset(btb_data_with_block_ram_1_reset),
    .io_wen(btb_data_with_block_ram_1_io_wen),
    .io_raddr(btb_data_with_block_ram_1_io_raddr),
    .io_waddr(btb_data_with_block_ram_1_io_waddr),
    .io_wdata(btb_data_with_block_ram_1_io_wdata),
    .io_rdata(btb_data_with_block_ram_1_io_rdata)
  );
  btb_data_with_block_ram btb_data_with_block_ram_2 ( // @[BTB.scala 250:54]
    .clock(btb_data_with_block_ram_2_clock),
    .reset(btb_data_with_block_ram_2_reset),
    .io_wen(btb_data_with_block_ram_2_io_wen),
    .io_raddr(btb_data_with_block_ram_2_io_raddr),
    .io_waddr(btb_data_with_block_ram_2_io_waddr),
    .io_wdata(btb_data_with_block_ram_2_io_wdata),
    .io_rdata(btb_data_with_block_ram_2_io_rdata)
  );
  btb_data_with_block_ram btb_data_with_block_ram_3 ( // @[BTB.scala 250:54]
    .clock(btb_data_with_block_ram_3_clock),
    .reset(btb_data_with_block_ram_3_reset),
    .io_wen(btb_data_with_block_ram_3_io_wen),
    .io_raddr(btb_data_with_block_ram_3_io_raddr),
    .io_waddr(btb_data_with_block_ram_3_io_waddr),
    .io_wdata(btb_data_with_block_ram_3_io_wdata),
    .io_rdata(btb_data_with_block_ram_3_io_rdata)
  );
  assign io_out_L = 2'h3 == ar_addr_reg[3:2] ? btb_banks_3_rdata : _GEN_2; // @[BTB.scala 265:{14,14}]
  assign io_hit_L = _GEN_15[3:0] == io_ar_addr_L[16:13] & _GEN_15[4]; // @[BTB.scala 286:167]
  assign btb_tag_with_block_ram_clock = clock;
  assign btb_tag_with_block_ram_reset = reset;
  assign btb_tag_with_block_ram_io_wen = _btb_banks_0_wen_T_1 & io_write; // @[BTB.scala 271:75]
  assign btb_tag_with_block_ram_io_raddr = io_ar_addr_L[12:4]; // @[BTB.scala 273:43]
  assign btb_tag_with_block_ram_io_waddr = io_aw_addr[12:4]; // @[BTB.scala 279:41]
  assign btb_tag_with_block_ram_io_wdata = {{3'd0}, _tag_banks_0_wdata_T_1}; // @[BTB.scala 249:28 272:28]
  assign btb_tag_with_block_ram_1_clock = clock;
  assign btb_tag_with_block_ram_1_reset = reset;
  assign btb_tag_with_block_ram_1_io_wen = _btb_banks_1_wen_T_1 & io_write; // @[BTB.scala 271:75]
  assign btb_tag_with_block_ram_1_io_raddr = io_ar_addr_L[12:4]; // @[BTB.scala 273:43]
  assign btb_tag_with_block_ram_1_io_waddr = io_aw_addr[12:4]; // @[BTB.scala 279:41]
  assign btb_tag_with_block_ram_1_io_wdata = {{3'd0}, _tag_banks_0_wdata_T_1}; // @[BTB.scala 249:28 272:28]
  assign btb_tag_with_block_ram_2_clock = clock;
  assign btb_tag_with_block_ram_2_reset = reset;
  assign btb_tag_with_block_ram_2_io_wen = _btb_banks_2_wen_T_1 & io_write; // @[BTB.scala 271:75]
  assign btb_tag_with_block_ram_2_io_raddr = io_ar_addr_L[12:4]; // @[BTB.scala 273:43]
  assign btb_tag_with_block_ram_2_io_waddr = io_aw_addr[12:4]; // @[BTB.scala 279:41]
  assign btb_tag_with_block_ram_2_io_wdata = {{3'd0}, _tag_banks_0_wdata_T_1}; // @[BTB.scala 249:28 272:28]
  assign btb_tag_with_block_ram_3_clock = clock;
  assign btb_tag_with_block_ram_3_reset = reset;
  assign btb_tag_with_block_ram_3_io_wen = _btb_banks_3_wen_T_1 & io_write; // @[BTB.scala 271:75]
  assign btb_tag_with_block_ram_3_io_raddr = io_ar_addr_L[12:4]; // @[BTB.scala 273:43]
  assign btb_tag_with_block_ram_3_io_waddr = io_aw_addr[12:4]; // @[BTB.scala 279:41]
  assign btb_tag_with_block_ram_3_io_wdata = {{3'd0}, _tag_banks_0_wdata_T_1}; // @[BTB.scala 249:28 272:28]
  assign btb_data_with_block_ram_clock = clock;
  assign btb_data_with_block_ram_reset = reset;
  assign btb_data_with_block_ram_io_wen = io_aw_addr[3:2] == 2'h0 & io_write; // @[BTB.scala 253:75]
  assign btb_data_with_block_ram_io_raddr = io_ar_addr_L[12:4]; // @[BTB.scala 255:43]
  assign btb_data_with_block_ram_io_waddr = io_aw_addr[12:4]; // @[BTB.scala 261:41]
  assign btb_data_with_block_ram_io_wdata = io_aw_target_addr; // @[BTB.scala 250:28 254:28]
  assign btb_data_with_block_ram_1_clock = clock;
  assign btb_data_with_block_ram_1_reset = reset;
  assign btb_data_with_block_ram_1_io_wen = io_aw_addr[3:2] == 2'h1 & io_write; // @[BTB.scala 253:75]
  assign btb_data_with_block_ram_1_io_raddr = io_ar_addr_L[12:4]; // @[BTB.scala 255:43]
  assign btb_data_with_block_ram_1_io_waddr = io_aw_addr[12:4]; // @[BTB.scala 261:41]
  assign btb_data_with_block_ram_1_io_wdata = io_aw_target_addr; // @[BTB.scala 250:28 254:28]
  assign btb_data_with_block_ram_2_clock = clock;
  assign btb_data_with_block_ram_2_reset = reset;
  assign btb_data_with_block_ram_2_io_wen = io_aw_addr[3:2] == 2'h2 & io_write; // @[BTB.scala 253:75]
  assign btb_data_with_block_ram_2_io_raddr = io_ar_addr_L[12:4]; // @[BTB.scala 255:43]
  assign btb_data_with_block_ram_2_io_waddr = io_aw_addr[12:4]; // @[BTB.scala 261:41]
  assign btb_data_with_block_ram_2_io_wdata = io_aw_target_addr; // @[BTB.scala 250:28 254:28]
  assign btb_data_with_block_ram_3_clock = clock;
  assign btb_data_with_block_ram_3_reset = reset;
  assign btb_data_with_block_ram_3_io_wen = io_aw_addr[3:2] == 2'h3 & io_write; // @[BTB.scala 253:75]
  assign btb_data_with_block_ram_3_io_raddr = io_ar_addr_L[12:4]; // @[BTB.scala 255:43]
  assign btb_data_with_block_ram_3_io_waddr = io_aw_addr[12:4]; // @[BTB.scala 261:41]
  assign btb_data_with_block_ram_3_io_wdata = io_aw_target_addr; // @[BTB.scala 250:28 254:28]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[BTB.scala 263:30]
      ar_addr_reg <= 64'h0; // @[BTB.scala 263:30]
    end else begin
      ar_addr_reg <= io_ar_addr_L; // @[BTB.scala 264:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  ar_addr_reg = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    ar_addr_reg = 64'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module branch_prediction_with_blockram(
  input         clock,
  input         reset,
  input  [63:0] io_pc,
  input  [63:0] io_write_pc,
  input  [3:0]  io_aw_pht_ways_addr,
  input  [6:0]  io_aw_pht_addr,
  input  [6:0]  io_aw_bht_addr,
  input  [63:0] io_aw_target_addr,
  input         io_btb_write,
  input         io_bht_write,
  input         io_pht_write,
  input  [6:0]  io_bht_in,
  input  [7:0]  io_pht_in,
  output [1:0]  io_out_L,
  output        io_pre_L,
  output [6:0]  io_bht_L,
  output        io_btb_hit_0,
  output [63:0] io_pre_target_L,
  input         io_stage2_stall,
  input         io_stage2_flush,
  output [7:0]  io_pht_lookup_value_out,
  output [6:0]  io_lookup_data_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  PHTS_banks_oneissue_block_ram_clock; // @[branch_prediction.scala 200:28]
  wire  PHTS_banks_oneissue_block_ram_reset; // @[branch_prediction.scala 200:28]
  wire [1:0] PHTS_banks_oneissue_block_ram_io_ar_bank_sel; // @[branch_prediction.scala 200:28]
  wire [6:0] PHTS_banks_oneissue_block_ram_io_ar_addr_L; // @[branch_prediction.scala 200:28]
  wire [2:0] PHTS_banks_oneissue_block_ram_io_ar_pht_addr; // @[branch_prediction.scala 200:28]
  wire [6:0] PHTS_banks_oneissue_block_ram_io_aw_addr; // @[branch_prediction.scala 200:28]
  wire [2:0] PHTS_banks_oneissue_block_ram_io_aw_pht_addr; // @[branch_prediction.scala 200:28]
  wire [1:0] PHTS_banks_oneissue_block_ram_io_aw_bank_sel; // @[branch_prediction.scala 200:28]
  wire  PHTS_banks_oneissue_block_ram_io_write; // @[branch_prediction.scala 200:28]
  wire [7:0] PHTS_banks_oneissue_block_ram_io_in; // @[branch_prediction.scala 200:28]
  wire [1:0] PHTS_banks_oneissue_block_ram_io_out_L; // @[branch_prediction.scala 200:28]
  wire [7:0] PHTS_banks_oneissue_block_ram_io_pht_out; // @[branch_prediction.scala 200:28]
  wire  BHT_banks_oneissue_clock; // @[branch_prediction.scala 201:28]
  wire  BHT_banks_oneissue_reset; // @[branch_prediction.scala 201:28]
  wire [1:0] BHT_banks_oneissue_io_ar_bank_sel; // @[branch_prediction.scala 201:28]
  wire [6:0] BHT_banks_oneissue_io_ar_addr_L; // @[branch_prediction.scala 201:28]
  wire [6:0] BHT_banks_oneissue_io_aw_addr; // @[branch_prediction.scala 201:28]
  wire  BHT_banks_oneissue_io_write; // @[branch_prediction.scala 201:28]
  wire [2:0] BHT_banks_oneissue_io_in; // @[branch_prediction.scala 201:28]
  wire [2:0] BHT_banks_oneissue_io_out_L; // @[branch_prediction.scala 201:28]
  wire  BTB_banks_oneissue_with_block_ram_clock; // @[branch_prediction.scala 202:27]
  wire  BTB_banks_oneissue_with_block_ram_reset; // @[branch_prediction.scala 202:27]
  wire [63:0] BTB_banks_oneissue_with_block_ram_io_ar_addr_L; // @[branch_prediction.scala 202:27]
  wire [63:0] BTB_banks_oneissue_with_block_ram_io_aw_addr; // @[branch_prediction.scala 202:27]
  wire [63:0] BTB_banks_oneissue_with_block_ram_io_aw_target_addr; // @[branch_prediction.scala 202:27]
  wire  BTB_banks_oneissue_with_block_ram_io_write; // @[branch_prediction.scala 202:27]
  wire [63:0] BTB_banks_oneissue_with_block_ram_io_out_L; // @[branch_prediction.scala 202:27]
  wire  BTB_banks_oneissue_with_block_ram_io_hit_L; // @[branch_prediction.scala 202:27]
  wire  pc_hash_num_array_0 = ^io_pc[7:4]; // @[macros.scala 447:45]
  wire  pc_hash_num_array_1 = ^io_pc[11:8]; // @[macros.scala 447:45]
  wire  pc_hash_num_array_2 = ^io_pc[15:12]; // @[macros.scala 447:45]
  wire  pc_hash_num_array_3 = ^io_pc[19:16]; // @[macros.scala 447:45]
  wire [3:0] pc_hash = {pc_hash_num_array_3,pc_hash_num_array_2,pc_hash_num_array_1,pc_hash_num_array_0}; // @[macros.scala 449:13]
  reg [6:0] stage_2_pht_lookup_0; // @[branch_prediction.scala 204:37]
  wire [6:0] stage_1_pht_lookup_0 = {BHT_banks_oneissue_io_out_L,io_pc[14:11]}; // @[Cat.scala 31:58]
  wire  _io_pre_L_T_1 = 2'h0 == io_out_L ? 1'h0 : 1'h1; // @[Mux.scala 81:58]
  wire  _io_pre_L_T_3 = 2'h1 == io_out_L ? 1'h0 : _io_pre_L_T_1; // @[Mux.scala 81:58]
  PHTS_banks_oneissue_block_ram PHTS_banks_oneissue_block_ram ( // @[branch_prediction.scala 200:28]
    .clock(PHTS_banks_oneissue_block_ram_clock),
    .reset(PHTS_banks_oneissue_block_ram_reset),
    .io_ar_bank_sel(PHTS_banks_oneissue_block_ram_io_ar_bank_sel),
    .io_ar_addr_L(PHTS_banks_oneissue_block_ram_io_ar_addr_L),
    .io_ar_pht_addr(PHTS_banks_oneissue_block_ram_io_ar_pht_addr),
    .io_aw_addr(PHTS_banks_oneissue_block_ram_io_aw_addr),
    .io_aw_pht_addr(PHTS_banks_oneissue_block_ram_io_aw_pht_addr),
    .io_aw_bank_sel(PHTS_banks_oneissue_block_ram_io_aw_bank_sel),
    .io_write(PHTS_banks_oneissue_block_ram_io_write),
    .io_in(PHTS_banks_oneissue_block_ram_io_in),
    .io_out_L(PHTS_banks_oneissue_block_ram_io_out_L),
    .io_pht_out(PHTS_banks_oneissue_block_ram_io_pht_out)
  );
  BHT_banks_oneissue BHT_banks_oneissue ( // @[branch_prediction.scala 201:28]
    .clock(BHT_banks_oneissue_clock),
    .reset(BHT_banks_oneissue_reset),
    .io_ar_bank_sel(BHT_banks_oneissue_io_ar_bank_sel),
    .io_ar_addr_L(BHT_banks_oneissue_io_ar_addr_L),
    .io_aw_addr(BHT_banks_oneissue_io_aw_addr),
    .io_write(BHT_banks_oneissue_io_write),
    .io_in(BHT_banks_oneissue_io_in),
    .io_out_L(BHT_banks_oneissue_io_out_L)
  );
  BTB_banks_oneissue_with_block_ram BTB_banks_oneissue_with_block_ram ( // @[branch_prediction.scala 202:27]
    .clock(BTB_banks_oneissue_with_block_ram_clock),
    .reset(BTB_banks_oneissue_with_block_ram_reset),
    .io_ar_addr_L(BTB_banks_oneissue_with_block_ram_io_ar_addr_L),
    .io_aw_addr(BTB_banks_oneissue_with_block_ram_io_aw_addr),
    .io_aw_target_addr(BTB_banks_oneissue_with_block_ram_io_aw_target_addr),
    .io_write(BTB_banks_oneissue_with_block_ram_io_write),
    .io_out_L(BTB_banks_oneissue_with_block_ram_io_out_L),
    .io_hit_L(BTB_banks_oneissue_with_block_ram_io_hit_L)
  );
  assign io_out_L = PHTS_banks_oneissue_block_ram_io_out_L; // @[branch_prediction.scala 288:14]
  assign io_pre_L = 2'h2 == io_out_L | _io_pre_L_T_3; // @[Mux.scala 81:58]
  assign io_bht_L = {{4'd0}, BHT_banks_oneissue_io_out_L}; // @[branch_prediction.scala 292:14]
  assign io_btb_hit_0 = BTB_banks_oneissue_with_block_ram_io_hit_L; // @[branch_prediction.scala 304:19]
  assign io_pre_target_L = BTB_banks_oneissue_with_block_ram_io_out_L; // @[branch_prediction.scala 300:21]
  assign io_pht_lookup_value_out = PHTS_banks_oneissue_block_ram_io_pht_out; // @[branch_prediction.scala 308:29]
  assign io_lookup_data_0 = stage_2_pht_lookup_0; // @[branch_prediction.scala 229:23]
  assign PHTS_banks_oneissue_block_ram_clock = clock;
  assign PHTS_banks_oneissue_block_ram_reset = reset;
  assign PHTS_banks_oneissue_block_ram_io_ar_bank_sel = io_pc[3:2]; // @[branch_prediction.scala 243:36]
  assign PHTS_banks_oneissue_block_ram_io_ar_addr_L = {BHT_banks_oneissue_io_out_L,io_pc[14:11]}; // @[Cat.scala 31:58]
  assign PHTS_banks_oneissue_block_ram_io_ar_pht_addr = pc_hash[2:0]; // @[branch_prediction.scala 244:28]
  assign PHTS_banks_oneissue_block_ram_io_aw_addr = io_aw_pht_addr; // @[branch_prediction.scala 259:24]
  assign PHTS_banks_oneissue_block_ram_io_aw_pht_addr = io_aw_pht_ways_addr[2:0]; // @[branch_prediction.scala 260:28]
  assign PHTS_banks_oneissue_block_ram_io_aw_bank_sel = io_write_pc[3:2]; // @[branch_prediction.scala 261:42]
  assign PHTS_banks_oneissue_block_ram_io_write = io_pht_write; // @[branch_prediction.scala 262:22]
  assign PHTS_banks_oneissue_block_ram_io_in = io_pht_in; // @[branch_prediction.scala 263:19]
  assign BHT_banks_oneissue_clock = clock;
  assign BHT_banks_oneissue_reset = reset;
  assign BHT_banks_oneissue_io_ar_bank_sel = io_pc[3:2]; // @[branch_prediction.scala 235:36]
  assign BHT_banks_oneissue_io_ar_addr_L = io_pc[10:4]; // @[branch_prediction.scala 237:34]
  assign BHT_banks_oneissue_io_aw_addr = io_aw_bht_addr; // @[branch_prediction.scala 241:24]
  assign BHT_banks_oneissue_io_write = io_bht_write; // @[branch_prediction.scala 236:22]
  assign BHT_banks_oneissue_io_in = io_bht_in[2:0]; // @[branch_prediction.scala 240:19]
  assign BTB_banks_oneissue_with_block_ram_clock = clock;
  assign BTB_banks_oneissue_with_block_ram_reset = reset;
  assign BTB_banks_oneissue_with_block_ram_io_ar_addr_L = io_pc; // @[branch_prediction.scala 266:25]
  assign BTB_banks_oneissue_with_block_ram_io_aw_addr = io_write_pc; // @[branch_prediction.scala 269:25]
  assign BTB_banks_oneissue_with_block_ram_io_aw_target_addr = io_aw_target_addr; // @[branch_prediction.scala 270:30]
  assign BTB_banks_oneissue_with_block_ram_io_write = io_btb_write; // @[branch_prediction.scala 271:21]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[branch_prediction.scala 218:33]
      stage_2_pht_lookup_0 <= 7'h0;
    end else if (io_stage2_flush) begin // @[branch_prediction.scala 218:57]
      stage_2_pht_lookup_0 <= 7'h0;
    end else if (io_stage2_stall) begin
      stage_2_pht_lookup_0 <= stage_1_pht_lookup_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stage_2_pht_lookup_0 = _RAND_0[6:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    stage_2_pht_lookup_0 = 7'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module bru_detail(
  input         clock,
  input         reset,
  input         io_stall,
  input         io_flush,
  input  [1:0]  io_in_pht,
  input  [6:0]  io_in_bht,
  input  [3:0]  io_in_hashcode,
  input  [63:0] io_in_target_pc,
  input  [6:0]  io_in_lookup_data,
  input  [7:0]  io_in_pht_lookup_value,
  output [1:0]  io_out_pht,
  output [6:0]  io_out_bht,
  output [3:0]  io_out_hashcode,
  output [63:0] io_out_target_pc,
  output [6:0]  io_out_lookup_data,
  output [7:0]  io_out_pht_lookup_value
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] pht_value; // @[myCPU.scala 660:34]
  reg [6:0] bht_value; // @[myCPU.scala 661:34]
  reg [3:0] hashcode_value; // @[myCPU.scala 662:39]
  reg [63:0] target_pc_value; // @[myCPU.scala 663:40]
  reg [6:0] lookup_data_value; // @[myCPU.scala 664:42]
  reg [7:0] pht_lookup_value_data; // @[myCPU.scala 665:46]
  assign io_out_pht = pht_value; // @[myCPU.scala 674:20]
  assign io_out_bht = bht_value; // @[myCPU.scala 675:20]
  assign io_out_hashcode = hashcode_value; // @[myCPU.scala 676:25]
  assign io_out_target_pc = target_pc_value; // @[myCPU.scala 677:26]
  assign io_out_lookup_data = lookup_data_value; // @[myCPU.scala 678:28]
  assign io_out_pht_lookup_value = pht_lookup_value_data; // @[myCPU.scala 679:33]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[myCPU.scala 666:25]
      pht_value <= 2'h0;
    end else if (io_flush) begin // @[myCPU.scala 666:42]
      pht_value <= 2'h0;
    end else if (io_stall) begin
      pht_value <= io_in_pht;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[myCPU.scala 667:25]
      bht_value <= 7'h0;
    end else if (io_flush) begin // @[myCPU.scala 667:42]
      bht_value <= 7'h0;
    end else if (io_stall) begin
      bht_value <= io_in_bht;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[myCPU.scala 668:30]
      hashcode_value <= 4'h0;
    end else if (io_flush) begin // @[myCPU.scala 668:47]
      hashcode_value <= 4'h0;
    end else if (io_stall) begin
      hashcode_value <= io_in_hashcode;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[myCPU.scala 669:31]
      target_pc_value <= 64'h0;
    end else if (io_flush) begin // @[myCPU.scala 669:48]
      target_pc_value <= 64'h0;
    end else if (io_stall) begin
      target_pc_value <= io_in_target_pc;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[myCPU.scala 670:33]
      lookup_data_value <= 7'h0;
    end else if (io_flush) begin // @[myCPU.scala 670:50]
      lookup_data_value <= 7'h0;
    end else if (io_stall) begin
      lookup_data_value <= io_in_lookup_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[myCPU.scala 671:37]
      pht_lookup_value_data <= 8'h0;
    end else if (io_flush) begin // @[myCPU.scala 671:54]
      pht_lookup_value_data <= 8'h0;
    end else if (io_stall) begin
      pht_lookup_value_data <= io_in_pht_lookup_value;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pht_value = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  bht_value = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  hashcode_value = _RAND_2[3:0];
  _RAND_3 = {2{`RANDOM}};
  target_pc_value = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  lookup_data_value = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  pht_lookup_value_data = _RAND_5[7:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    pht_value = 2'h0;
  end
  if (reset) begin
    bht_value = 7'h0;
  end
  if (reset) begin
    hashcode_value = 4'h0;
  end
  if (reset) begin
    target_pc_value = 64'h0;
  end
  if (reset) begin
    lookup_data_value = 7'h0;
  end
  if (reset) begin
    pht_lookup_value_data = 8'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module myCPU(
  input         ext_int_timer,
  input         resetn,
  input         clk,
  output        inst_cache,
  output        inst_sram_en,
  output [63:0] inst_sram_addr,
  input  [39:0] inst_sram_rdata_L,
  input  [1:0]  inst_write_en,
  output        stage2_flush,
  input         stage2_stall,
  output        stage1_valid_flush,
  output        inst_ready_to_use,
  output        inst_buffer_full,
  output        data_sram_en,
  output        data_sram_wen,
  output [1:0]  data_size,
  output [63:0] data_sram_addr,
  output [63:0] data_sram_wdata,
  output        data_cache,
  input  [63:0] data_sram_rdata,
  input         data_stage2_stall,
  output [7:0]  data_wstrb,
  output        data_fence_i_control,
  output [63:0] debug_wb_pc,
  output [3:0]  debug_wb_rf_wen,
  output [4:0]  debug_wb_rf_wnum,
  output [63:0] debug_wb_rf_wdata,
  output        icache_tag_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [63:0] _RAND_36;
`endif // RANDOMIZE_REG_INIT
  wire [23:0] _alu_io_ctrl; // @[myCPU.scala 120:22]
  wire [63:0] _alu_io_in1; // @[myCPU.scala 120:22]
  wire [63:0] _alu_io_in2; // @[myCPU.scala 120:22]
  wire [63:0] _alu_io_result; // @[myCPU.scala 120:22]
  wire  _alu_io_overflow; // @[myCPU.scala 120:22]
  wire  _alu_io_data_w; // @[myCPU.scala 120:22]
  wire  _br_reset; // @[myCPU.scala 121:22]
  wire [63:0] _br_io_r1; // @[myCPU.scala 121:22]
  wire [63:0] _br_io_r2; // @[myCPU.scala 121:22]
  wire [5:0] _br_io_branch; // @[myCPU.scala 121:22]
  wire  _br_io_exe; // @[myCPU.scala 121:22]
  wire  _cfu_reset; // @[myCPU.scala 122:22]
  wire  _cfu_io_Inst_Fifo_Empty; // @[myCPU.scala 122:22]
  wire  _cfu_io_dmem_calD; // @[myCPU.scala 122:22]
  wire  _cfu_io_BranchD_Flag; // @[myCPU.scala 122:22]
  wire  _cfu_io_JRD; // @[myCPU.scala 122:22]
  wire  _cfu_io_CanBranchD; // @[myCPU.scala 122:22]
  wire  _cfu_io_DivPendingE; // @[myCPU.scala 122:22]
  wire  _cfu_io_DataPendingM; // @[myCPU.scala 122:22]
  wire  _cfu_io_InException; // @[myCPU.scala 122:22]
  wire [4:0] _cfu_io_WriteRegE; // @[myCPU.scala 122:22]
  wire  _cfu_io_RegWriteE; // @[myCPU.scala 122:22]
  wire  _cfu_io_csrToRegE; // @[myCPU.scala 122:22]
  wire [4:0] _cfu_io_WriteRegM; // @[myCPU.scala 122:22]
  wire  _cfu_io_MemToRegM; // @[myCPU.scala 122:22]
  wire  _cfu_io_RegWriteM; // @[myCPU.scala 122:22]
  wire  _cfu_io_csrWriteM; // @[myCPU.scala 122:22]
  wire [4:0] _cfu_io_WriteRegM2; // @[myCPU.scala 122:22]
  wire  _cfu_io_MemToRegM2; // @[myCPU.scala 122:22]
  wire  _cfu_io_RegWriteM2; // @[myCPU.scala 122:22]
  wire  _cfu_io_csrWriteM2; // @[myCPU.scala 122:22]
  wire [4:0] _cfu_io_WriteRegW; // @[myCPU.scala 122:22]
  wire  _cfu_io_RegWriteW; // @[myCPU.scala 122:22]
  wire [11:0] _cfu_io_ReadcsrAddrE; // @[myCPU.scala 122:22]
  wire [11:0] _cfu_io_WritecsrAddrM; // @[myCPU.scala 122:22]
  wire [11:0] _cfu_io_WritecsrAddrM2; // @[myCPU.scala 122:22]
  wire [4:0] _cfu_io_R2D; // @[myCPU.scala 122:22]
  wire [4:0] _cfu_io_R1D; // @[myCPU.scala 122:22]
  wire [4:0] _cfu_io_R2E; // @[myCPU.scala 122:22]
  wire [4:0] _cfu_io_R1E; // @[myCPU.scala 122:22]
  wire  _cfu_io_StallF; // @[myCPU.scala 122:22]
  wire  _cfu_io_StallD; // @[myCPU.scala 122:22]
  wire  _cfu_io_StallE; // @[myCPU.scala 122:22]
  wire  _cfu_io_StallM; // @[myCPU.scala 122:22]
  wire  _cfu_io_StallM2; // @[myCPU.scala 122:22]
  wire  _cfu_io_StallW; // @[myCPU.scala 122:22]
  wire  _cfu_io_FlushD; // @[myCPU.scala 122:22]
  wire  _cfu_io_FlushE; // @[myCPU.scala 122:22]
  wire  _cfu_io_FlushM; // @[myCPU.scala 122:22]
  wire  _cfu_io_FlushM2; // @[myCPU.scala 122:22]
  wire  _cfu_io_FlushW; // @[myCPU.scala 122:22]
  wire [1:0] _cfu_io_Forward1E; // @[myCPU.scala 122:22]
  wire [1:0] _cfu_io_Forward2E; // @[myCPU.scala 122:22]
  wire [1:0] _cfu_io_Forward1D; // @[myCPU.scala 122:22]
  wire [1:0] _cfu_io_Forward2D; // @[myCPU.scala 122:22]
  wire [1:0] _cfu_io_ForwardcsrE; // @[myCPU.scala 122:22]
  wire  _csr_clock; // @[myCPU.scala 123:22]
  wire  _csr_reset; // @[myCPU.scala 123:22]
  wire [11:0] _csr_io_csr_read_addr; // @[myCPU.scala 123:22]
  wire [11:0] _csr_io_csr_write_addr; // @[myCPU.scala 123:22]
  wire [63:0] _csr_io_csr_write_data; // @[myCPU.scala 123:22]
  wire  _csr_io_csr_write_en; // @[myCPU.scala 123:22]
  wire [63:0] _csr_io_pc; // @[myCPU.scala 123:22]
  wire [31:0] _csr_io_exception_type_i; // @[myCPU.scala 123:22]
  wire [63:0] _csr_io_return_pc; // @[myCPU.scala 123:22]
  wire  _csr_io_exception; // @[myCPU.scala 123:22]
  wire [63:0] _csr_io_csr_read_data; // @[myCPU.scala 123:22]
  wire  _csr_io_icache_tags_flush; // @[myCPU.scala 123:22]
  wire  _csr_io_int_type_timer; // @[myCPU.scala 123:22]
  wire  _csr_io_Int_able; // @[myCPU.scala 123:22]
  wire  _csr_io_int_type_able_timer; // @[myCPU.scala 123:22]
  wire [31:0] _cu_io1_InstrD; // @[myCPU.scala 124:22]
  wire  _cu_io1_BadInstrD; // @[myCPU.scala 124:22]
  wire  _cu_io1_SysCallD; // @[myCPU.scala 124:22]
  wire  _cu_io1_EretD; // @[myCPU.scala 124:22]
  wire  _cu_io1_dmem_addr_cal; // @[myCPU.scala 124:22]
  wire  _cu_io_RegWriteD; // @[myCPU.scala 124:22]
  wire  _cu_io_MemToRegD; // @[myCPU.scala 124:22]
  wire  _cu_io_MemWriteD; // @[myCPU.scala 124:22]
  wire [23:0] _cu_io_ALUCtrlD; // @[myCPU.scala 124:22]
  wire [1:0] _cu_io_ALUSrcD_0; // @[myCPU.scala 124:22]
  wire [1:0] _cu_io_ALUSrcD_1; // @[myCPU.scala 124:22]
  wire [4:0] _cu_io_RegDstD; // @[myCPU.scala 124:22]
  wire  _cu_io_LinkD; // @[myCPU.scala 124:22]
  wire  _cu_io_csrWriteD; // @[myCPU.scala 124:22]
  wire  _cu_io_csrToRegD; // @[myCPU.scala 124:22]
  wire  _cu_io_LoadUnsignedD; // @[myCPU.scala 124:22]
  wire [1:0] _cu_io_MemWidthD; // @[myCPU.scala 124:22]
  wire [63:0] _cu_io_ImmD; // @[myCPU.scala 124:22]
  wire  _cu_io_ebreakD; // @[myCPU.scala 124:22]
  wire  _cu_io_data_wD; // @[myCPU.scala 124:22]
  wire [23:0] _cu_io_muldiv_control; // @[myCPU.scala 124:22]
  wire  _cu_io_muldiv_cal; // @[myCPU.scala 124:22]
  wire  _cu_io_alu_cal; // @[myCPU.scala 124:22]
  wire [5:0] _cu_io_csr_control; // @[myCPU.scala 124:22]
  wire  _cu_io_csr_Imm; // @[myCPU.scala 124:22]
  wire  _cu_io_fence_i_control; // @[myCPU.scala 124:22]
  wire  _dmem_io_data_ok; // @[myCPU.scala 125:23]
  wire [63:0] _dmem_io_rdata; // @[myCPU.scala 125:23]
  wire [63:0] _dmem_io_Physisc_Address; // @[myCPU.scala 125:23]
  wire [1:0] _dmem_io_WIDTH; // @[myCPU.scala 125:23]
  wire  _dmem_io_SIGN; // @[myCPU.scala 125:23]
  wire [63:0] _dmem_io_RD; // @[myCPU.scala 125:23]
  wire  _dmem_io_data_pending; // @[myCPU.scala 125:23]
  wire  _dmemreq_io_en; // @[myCPU.scala 126:26]
  wire  _dmemreq_io_MemWriteE; // @[myCPU.scala 126:26]
  wire  _dmemreq_io_MemToRegE; // @[myCPU.scala 126:26]
  wire [1:0] _dmemreq_io_MemWidthE; // @[myCPU.scala 126:26]
  wire [63:0] _dmemreq_io_VAddrE; // @[myCPU.scala 126:26]
  wire [63:0] _dmemreq_io_WriteDataE; // @[myCPU.scala 126:26]
  wire  _dmemreq_io_req; // @[myCPU.scala 126:26]
  wire  _dmemreq_io_wr; // @[myCPU.scala 126:26]
  wire [1:0] _dmemreq_io_size; // @[myCPU.scala 126:26]
  wire [63:0] _dmemreq_io_addr; // @[myCPU.scala 126:26]
  wire [63:0] _dmemreq_io_wdata; // @[myCPU.scala 126:26]
  wire [7:0] _dmemreq_io_wstrb; // @[myCPU.scala 126:26]
  wire  _ex2mem_clock; // @[myCPU.scala 127:26]
  wire  _ex2mem_reset; // @[myCPU.scala 127:26]
  wire  _ex2mem_io1_RegWriteE; // @[myCPU.scala 127:26]
  wire  _ex2mem_io1_MemToRegE; // @[myCPU.scala 127:26]
  wire  _ex2mem_io1_LoadUnsignedE; // @[myCPU.scala 127:26]
  wire [1:0] _ex2mem_io1_MemWidthE; // @[myCPU.scala 127:26]
  wire  _ex2mem_io1_csrWriteE; // @[myCPU.scala 127:26]
  wire [11:0] _ex2mem_io1_WritecsrAddrE; // @[myCPU.scala 127:26]
  wire [63:0] _ex2mem_io1_PCE; // @[myCPU.scala 127:26]
  wire [1:0] _ex2mem_io1_MemRLE; // @[myCPU.scala 127:26]
  wire [1:0] _ex2mem_io1_BranchJump_JrE; // @[myCPU.scala 127:26]
  wire [2:0] _ex2mem_io1_Tlb_Control; // @[myCPU.scala 127:26]
  wire  _ex2mem_io1_eBreakE; // @[myCPU.scala 127:26]
  wire  _ex2mem_io1_fence_i_control; // @[myCPU.scala 127:26]
  wire  _ex2mem_io_en; // @[myCPU.scala 127:26]
  wire  _ex2mem_io_clr; // @[myCPU.scala 127:26]
  wire [63:0] _ex2mem_io_WriteDataE; // @[myCPU.scala 127:26]
  wire [4:0] _ex2mem_io_WriteRegE; // @[myCPU.scala 127:26]
  wire [63:0] _ex2mem_io_PhyAddrE; // @[myCPU.scala 127:26]
  wire [63:0] _ex2mem_io_CsrWritedataE; // @[myCPU.scala 127:26]
  wire [31:0] _ex2mem_io_ExceptionTypeE; // @[myCPU.scala 127:26]
  wire [63:0] _ex2mem_io_RtE; // @[myCPU.scala 127:26]
  wire [63:0] _ex2mem_io_Pc_NextE; // @[myCPU.scala 127:26]
  wire [63:0] _ex2mem_io_mem_trace_budleE_pc; // @[myCPU.scala 127:26]
  wire [63:0] _ex2mem_io_mem_trace_budleE_data; // @[myCPU.scala 127:26]
  wire [1:0] _ex2mem_io_mem_trace_budleE_mem_fetch_type; // @[myCPU.scala 127:26]
  wire [63:0] _ex2mem_io_mem_trace_budleE_addr; // @[myCPU.scala 127:26]
  wire [2:0] _ex2mem_io_mem_trace_budleE_len; // @[myCPU.scala 127:26]
  wire  _ex2mem_io_mem_trace_budleE_cache; // @[myCPU.scala 127:26]
  wire  _ex2mem_io_RegWriteM; // @[myCPU.scala 127:26]
  wire  _ex2mem_io_MemToRegM; // @[myCPU.scala 127:26]
  wire [63:0] _ex2mem_io_WriteDataM; // @[myCPU.scala 127:26]
  wire [4:0] _ex2mem_io_WriteRegM; // @[myCPU.scala 127:26]
  wire  _ex2mem_io_LoadUnsignedM; // @[myCPU.scala 127:26]
  wire [1:0] _ex2mem_io_MemWidthM; // @[myCPU.scala 127:26]
  wire [63:0] _ex2mem_io_PhyAddrM; // @[myCPU.scala 127:26]
  wire  _ex2mem_io_csrWriteM; // @[myCPU.scala 127:26]
  wire [11:0] _ex2mem_io_WritecsrAddrM; // @[myCPU.scala 127:26]
  wire [63:0] _ex2mem_io_PCM; // @[myCPU.scala 127:26]
  wire [31:0] _ex2mem_io_ExceptionTypeM_Out; // @[myCPU.scala 127:26]
  wire [1:0] _ex2mem_io_MemRLM; // @[myCPU.scala 127:26]
  wire [63:0] _ex2mem_io_RtM; // @[myCPU.scala 127:26]
  wire [1:0] _ex2mem_io_BranchJump_JrM; // @[myCPU.scala 127:26]
  wire [2:0] _ex2mem_io_Tlb_ControlM; // @[myCPU.scala 127:26]
  wire  _ex2mem_io_eBreakM; // @[myCPU.scala 127:26]
  wire [63:0] _ex2mem_io_Pc_NextM; // @[myCPU.scala 127:26]
  wire [63:0] _ex2mem_io_mem_trace_budleM_pc; // @[myCPU.scala 127:26]
  wire [63:0] _ex2mem_io_mem_trace_budleM_data; // @[myCPU.scala 127:26]
  wire [1:0] _ex2mem_io_mem_trace_budleM_mem_fetch_type; // @[myCPU.scala 127:26]
  wire [63:0] _ex2mem_io_mem_trace_budleM_addr; // @[myCPU.scala 127:26]
  wire [2:0] _ex2mem_io_mem_trace_budleM_len; // @[myCPU.scala 127:26]
  wire  _ex2mem_io_mem_trace_budleM_cache; // @[myCPU.scala 127:26]
  wire [63:0] _ex2mem_io_CsrWritedataM; // @[myCPU.scala 127:26]
  wire  _ex2mem_io_fence_i_controlM; // @[myCPU.scala 127:26]
  wire  _mem2mem2_clock; // @[myCPU.scala 128:28]
  wire  _mem2mem2_reset; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io1_RegWriteE; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io1_MemToRegE; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io1_LoadUnsignedE; // @[myCPU.scala 128:28]
  wire [1:0] _mem2mem2_io1_MemWidthE; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io1_csrWriteE; // @[myCPU.scala 128:28]
  wire [11:0] _mem2mem2_io1_WritecsrAddrE; // @[myCPU.scala 128:28]
  wire [63:0] _mem2mem2_io1_PCE; // @[myCPU.scala 128:28]
  wire [1:0] _mem2mem2_io1_MemRLE; // @[myCPU.scala 128:28]
  wire [1:0] _mem2mem2_io1_BranchJump_JrE; // @[myCPU.scala 128:28]
  wire [2:0] _mem2mem2_io1_Tlb_Control; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io1_eBreakE; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io1_fence_i_control; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io_en; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io_clr; // @[myCPU.scala 128:28]
  wire [63:0] _mem2mem2_io_WriteDataE; // @[myCPU.scala 128:28]
  wire [4:0] _mem2mem2_io_WriteRegE; // @[myCPU.scala 128:28]
  wire [63:0] _mem2mem2_io_PhyAddrE; // @[myCPU.scala 128:28]
  wire [63:0] _mem2mem2_io_CsrWritedataE; // @[myCPU.scala 128:28]
  wire [31:0] _mem2mem2_io_ExceptionTypeE; // @[myCPU.scala 128:28]
  wire [63:0] _mem2mem2_io_RtE; // @[myCPU.scala 128:28]
  wire [63:0] _mem2mem2_io_Pc_NextE; // @[myCPU.scala 128:28]
  wire [63:0] _mem2mem2_io_mem_trace_budleE_pc; // @[myCPU.scala 128:28]
  wire [63:0] _mem2mem2_io_mem_trace_budleE_data; // @[myCPU.scala 128:28]
  wire [1:0] _mem2mem2_io_mem_trace_budleE_mem_fetch_type; // @[myCPU.scala 128:28]
  wire [63:0] _mem2mem2_io_mem_trace_budleE_addr; // @[myCPU.scala 128:28]
  wire [2:0] _mem2mem2_io_mem_trace_budleE_len; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io_mem_trace_budleE_cache; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io_RegWriteM; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io_MemToRegM; // @[myCPU.scala 128:28]
  wire [63:0] _mem2mem2_io_WriteDataM; // @[myCPU.scala 128:28]
  wire [4:0] _mem2mem2_io_WriteRegM; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io_LoadUnsignedM; // @[myCPU.scala 128:28]
  wire [1:0] _mem2mem2_io_MemWidthM; // @[myCPU.scala 128:28]
  wire [63:0] _mem2mem2_io_PhyAddrM; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io_csrWriteM; // @[myCPU.scala 128:28]
  wire [11:0] _mem2mem2_io_WritecsrAddrM; // @[myCPU.scala 128:28]
  wire [63:0] _mem2mem2_io_PCM; // @[myCPU.scala 128:28]
  wire [31:0] _mem2mem2_io_ExceptionTypeM_Out; // @[myCPU.scala 128:28]
  wire [1:0] _mem2mem2_io_MemRLM; // @[myCPU.scala 128:28]
  wire [63:0] _mem2mem2_io_RtM; // @[myCPU.scala 128:28]
  wire [1:0] _mem2mem2_io_BranchJump_JrM; // @[myCPU.scala 128:28]
  wire [2:0] _mem2mem2_io_Tlb_ControlM; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io_eBreakM; // @[myCPU.scala 128:28]
  wire [63:0] _mem2mem2_io_Pc_NextM; // @[myCPU.scala 128:28]
  wire [63:0] _mem2mem2_io_mem_trace_budleM_pc; // @[myCPU.scala 128:28]
  wire [63:0] _mem2mem2_io_mem_trace_budleM_data; // @[myCPU.scala 128:28]
  wire [1:0] _mem2mem2_io_mem_trace_budleM_mem_fetch_type; // @[myCPU.scala 128:28]
  wire [63:0] _mem2mem2_io_mem_trace_budleM_addr; // @[myCPU.scala 128:28]
  wire [2:0] _mem2mem2_io_mem_trace_budleM_len; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io_mem_trace_budleM_cache; // @[myCPU.scala 128:28]
  wire [63:0] _mem2mem2_io_CsrWritedataM; // @[myCPU.scala 128:28]
  wire  _mem2mem2_io_fence_i_controlM; // @[myCPU.scala 128:28]
  wire  _id2ex_clock; // @[myCPU.scala 130:26]
  wire  _id2ex_reset; // @[myCPU.scala 130:26]
  wire  _id2ex_io1_RegWriteD; // @[myCPU.scala 130:26]
  wire  _id2ex_io1_MemToRegD; // @[myCPU.scala 130:26]
  wire  _id2ex_io1_MemWriteD; // @[myCPU.scala 130:26]
  wire [23:0] _id2ex_io1_ALUCtrlD; // @[myCPU.scala 130:26]
  wire [1:0] _id2ex_io1_ALUSrcD_0; // @[myCPU.scala 130:26]
  wire [1:0] _id2ex_io1_ALUSrcD_1; // @[myCPU.scala 130:26]
  wire [4:0] _id2ex_io1_RegDstD; // @[myCPU.scala 130:26]
  wire  _id2ex_io1_LinkD; // @[myCPU.scala 130:26]
  wire  _id2ex_io1_csrWriteD; // @[myCPU.scala 130:26]
  wire  _id2ex_io1_csrToRegD; // @[myCPU.scala 130:26]
  wire  _id2ex_io1_LoadUnsignedD; // @[myCPU.scala 130:26]
  wire [1:0] _id2ex_io1_MemWidthD; // @[myCPU.scala 130:26]
  wire  _id2ex_io1_ebreakD; // @[myCPU.scala 130:26]
  wire  _id2ex_io1_data_wD; // @[myCPU.scala 130:26]
  wire [23:0] _id2ex_io1_muldiv_control; // @[myCPU.scala 130:26]
  wire  _id2ex_io1_muldiv_cal; // @[myCPU.scala 130:26]
  wire  _id2ex_io1_alu_cal; // @[myCPU.scala 130:26]
  wire [5:0] _id2ex_io1_csr_control; // @[myCPU.scala 130:26]
  wire  _id2ex_io1_csr_Imm; // @[myCPU.scala 130:26]
  wire  _id2ex_io1_fence_i_control; // @[myCPU.scala 130:26]
  wire  _id2ex_io2_RegWriteE; // @[myCPU.scala 130:26]
  wire  _id2ex_io2_MemToRegE; // @[myCPU.scala 130:26]
  wire  _id2ex_io2_MemWriteE; // @[myCPU.scala 130:26]
  wire [23:0] _id2ex_io2_ALUCtrlE; // @[myCPU.scala 130:26]
  wire  _id2ex_io2_ALUSrcE_0; // @[myCPU.scala 130:26]
  wire  _id2ex_io2_ALUSrcE_1; // @[myCPU.scala 130:26]
  wire [4:0] _id2ex_io2_RegDstE; // @[myCPU.scala 130:26]
  wire  _id2ex_io2_LinkE; // @[myCPU.scala 130:26]
  wire [63:0] _id2ex_io2_PCPlus4E; // @[myCPU.scala 130:26]
  wire  _id2ex_io2_LoadUnsignedE; // @[myCPU.scala 130:26]
  wire [1:0] _id2ex_io2_MemWidthE; // @[myCPU.scala 130:26]
  wire  _id2ex_io2_csrWriteE; // @[myCPU.scala 130:26]
  wire [11:0] _id2ex_io2_WritecsrAddrE; // @[myCPU.scala 130:26]
  wire [11:0] _id2ex_io2_ReadcsrAddrE; // @[myCPU.scala 130:26]
  wire [63:0] _id2ex_io2_PCE; // @[myCPU.scala 130:26]
  wire [1:0] _id2ex_io2_BranchJump_JrE; // @[myCPU.scala 130:26]
  wire  _id2ex_io2_eBreakE; // @[myCPU.scala 130:26]
  wire  _id2ex_io2_fence_i_control; // @[myCPU.scala 130:26]
  wire  _id2ex_io_en; // @[myCPU.scala 130:26]
  wire  _id2ex_io_clr; // @[myCPU.scala 130:26]
  wire  _id2ex_io_csrToRegE_Out; // @[myCPU.scala 130:26]
  wire [63:0] _id2ex_io_RD1D; // @[myCPU.scala 130:26]
  wire [63:0] _id2ex_io_RD2D; // @[myCPU.scala 130:26]
  wire [4:0] _id2ex_io_R2D; // @[myCPU.scala 130:26]
  wire [4:0] _id2ex_io_R1D; // @[myCPU.scala 130:26]
  wire [63:0] _id2ex_io_ImmD; // @[myCPU.scala 130:26]
  wire [63:0] _id2ex_io_PCPlus4D; // @[myCPU.scala 130:26]
  wire [11:0] _id2ex_io_WritecsrAddrD; // @[myCPU.scala 130:26]
  wire [11:0] _id2ex_io_ReadcsrAddrD; // @[myCPU.scala 130:26]
  wire [63:0] _id2ex_io_PCD; // @[myCPU.scala 130:26]
  wire [31:0] _id2ex_io_ExceptionTypeD; // @[myCPU.scala 130:26]
  wire [63:0] _id2ex_io_Pc_NextD; // @[myCPU.scala 130:26]
  wire [1:0] _id2ex_io_BranchJump_JrD; // @[myCPU.scala 130:26]
  wire [63:0] _id2ex_io_RD1E; // @[myCPU.scala 130:26]
  wire [63:0] _id2ex_io_RD2E; // @[myCPU.scala 130:26]
  wire [4:0] _id2ex_io_R2E; // @[myCPU.scala 130:26]
  wire [4:0] _id2ex_io_R1E; // @[myCPU.scala 130:26]
  wire [63:0] _id2ex_io_ImmE; // @[myCPU.scala 130:26]
  wire  _id2ex_io_data_wE; // @[myCPU.scala 130:26]
  wire [63:0] _id2ex_io_Pc_NextE; // @[myCPU.scala 130:26]
  wire [23:0] _id2ex_io_muldiv_control; // @[myCPU.scala 130:26]
  wire  _id2ex_io_alu_calE; // @[myCPU.scala 130:26]
  wire  _id2ex_io_muldiv_calE; // @[myCPU.scala 130:26]
  wire [31:0] _id2ex_io_ExceptionTypeE_Out; // @[myCPU.scala 130:26]
  wire [5:0] _id2ex_io_csr_controlE; // @[myCPU.scala 130:26]
  wire  _id2ex_io_csr_ImmE; // @[myCPU.scala 130:26]
  wire  _if2id_clock; // @[myCPU.scala 131:26]
  wire  _if2id_reset; // @[myCPU.scala 131:26]
  wire  _if2id_io_en; // @[myCPU.scala 131:26]
  wire  _if2id_io_clr; // @[myCPU.scala 131:26]
  wire [63:0] _if2id_io_InstrF; // @[myCPU.scala 131:26]
  wire [63:0] _if2id_io_PCPlus4F; // @[myCPU.scala 131:26]
  wire [63:0] _if2id_io_PCF; // @[myCPU.scala 131:26]
  wire [1:0] _if2id_io_ExceptionTypeF; // @[myCPU.scala 131:26]
  wire [31:0] _if2id_io_InstrD; // @[myCPU.scala 131:26]
  wire [63:0] _if2id_io_PCPlus4D; // @[myCPU.scala 131:26]
  wire [63:0] _if2id_io_PCD; // @[myCPU.scala 131:26]
  wire [1:0] _if2id_io_ExceptionTypeD_Out; // @[myCPU.scala 131:26]
  wire  _mem22wb_clock; // @[myCPU.scala 133:27]
  wire  _mem22wb_reset; // @[myCPU.scala 133:27]
  wire  _mem22wb_io_en; // @[myCPU.scala 133:27]
  wire  _mem22wb_io_clr; // @[myCPU.scala 133:27]
  wire  _mem22wb_io_RegWriteM; // @[myCPU.scala 133:27]
  wire [63:0] _mem22wb_io_ResultM; // @[myCPU.scala 133:27]
  wire [4:0] _mem22wb_io_WriteRegM; // @[myCPU.scala 133:27]
  wire  _mem22wb_io_csrWriteM; // @[myCPU.scala 133:27]
  wire [11:0] _mem22wb_io_WritecsrAddrM; // @[myCPU.scala 133:27]
  wire [63:0] _mem22wb_io_CsrWritedataM; // @[myCPU.scala 133:27]
  wire [63:0] _mem22wb_io_PCM; // @[myCPU.scala 133:27]
  wire [31:0] _mem22wb_io_ExceptionTypeM; // @[myCPU.scala 133:27]
  wire [1:0] _mem22wb_io_BranchJump_JrM; // @[myCPU.scala 133:27]
  wire  _mem22wb_io_eBreakM; // @[myCPU.scala 133:27]
  wire [63:0] _mem22wb_io_Pc_NextM; // @[myCPU.scala 133:27]
  wire [63:0] _mem22wb_io_Mem_trace_budleM_pc; // @[myCPU.scala 133:27]
  wire [63:0] _mem22wb_io_Mem_trace_budleM_data; // @[myCPU.scala 133:27]
  wire [1:0] _mem22wb_io_Mem_trace_budleM_mem_fetch_type; // @[myCPU.scala 133:27]
  wire [63:0] _mem22wb_io_Mem_trace_budleM_addr; // @[myCPU.scala 133:27]
  wire [2:0] _mem22wb_io_Mem_trace_budleM_len; // @[myCPU.scala 133:27]
  wire  _mem22wb_io_Mem_trace_budleM_cache; // @[myCPU.scala 133:27]
  wire  _mem22wb_io_RegWriteW_Out; // @[myCPU.scala 133:27]
  wire [63:0] _mem22wb_io_ResultW; // @[myCPU.scala 133:27]
  wire [4:0] _mem22wb_io_WriteRegW; // @[myCPU.scala 133:27]
  wire  _mem22wb_io_csrWriteW; // @[myCPU.scala 133:27]
  wire [11:0] _mem22wb_io_WritecsrAddrW; // @[myCPU.scala 133:27]
  wire [63:0] _mem22wb_io_PCW; // @[myCPU.scala 133:27]
  wire [31:0] _mem22wb_io_ExceptionTypeW_Out; // @[myCPU.scala 133:27]
  wire [1:0] _mem22wb_io_BranchJump_JrW; // @[myCPU.scala 133:27]
  wire  _mem22wb_io_eBreakW; // @[myCPU.scala 133:27]
  wire [63:0] _mem22wb_io_Pc_NextW; // @[myCPU.scala 133:27]
  wire [63:0] _mem22wb_io_Mem_trace_budleW_pc; // @[myCPU.scala 133:27]
  wire [63:0] _mem22wb_io_Mem_trace_budleW_data; // @[myCPU.scala 133:27]
  wire [1:0] _mem22wb_io_Mem_trace_budleW_mem_fetch_type; // @[myCPU.scala 133:27]
  wire [63:0] _mem22wb_io_Mem_trace_budleW_addr; // @[myCPU.scala 133:27]
  wire [2:0] _mem22wb_io_Mem_trace_budleW_len; // @[myCPU.scala 133:27]
  wire  _mem22wb_io_Mem_trace_budleW_cache; // @[myCPU.scala 133:27]
  wire [63:0] _mem22wb_io_CsrWritedataW; // @[myCPU.scala 133:27]
  wire [63:0] _addr_cal_io_d_vaddr; // @[myCPU.scala 134:31]
  wire [63:0] _addr_cal_io_d_paddr; // @[myCPU.scala 134:31]
  wire  _addr_cal_io_d_cached; // @[myCPU.scala 134:31]
  wire  _muldiv_clock; // @[myCPU.scala 135:26]
  wire  _muldiv_reset; // @[myCPU.scala 135:26]
  wire  _muldiv_io_en; // @[myCPU.scala 135:26]
  wire [23:0] _muldiv_io_ctrl; // @[myCPU.scala 135:26]
  wire [63:0] _muldiv_io_in1; // @[myCPU.scala 135:26]
  wire [63:0] _muldiv_io_in2; // @[myCPU.scala 135:26]
  wire [63:0] _muldiv_io_data_out; // @[myCPU.scala 135:26]
  wire  _muldiv_io_pending; // @[myCPU.scala 135:26]
  wire  _regfile_clock; // @[myCPU.scala 137:26]
  wire  _regfile_reset; // @[myCPU.scala 137:26]
  wire [4:0] _regfile_io_A1; // @[myCPU.scala 137:26]
  wire [4:0] _regfile_io_A2; // @[myCPU.scala 137:26]
  wire  _regfile_io_WE3; // @[myCPU.scala 137:26]
  wire [4:0] _regfile_io_A3; // @[myCPU.scala 137:26]
  wire [63:0] _regfile_io_WD3; // @[myCPU.scala 137:26]
  wire [63:0] _regfile_io_RD1; // @[myCPU.scala 137:26]
  wire [63:0] _regfile_io_RD2; // @[myCPU.scala 137:26]
  wire [2047:0] _regfile_io_reg_file_alL_out; // @[myCPU.scala 137:26]
  wire  _mtrace_mod_reset; // @[myCPU.scala 138:29]
  wire  _mtrace_mod_clock; // @[myCPU.scala 138:29]
  wire [63:0] _mtrace_mod_data; // @[myCPU.scala 138:29]
  wire [63:0] _mtrace_mod_pc; // @[myCPU.scala 138:29]
  wire [63:0] _mtrace_mod_addr; // @[myCPU.scala 138:29]
  wire  _mtrace_mod_mem_req; // @[myCPU.scala 138:29]
  wire  _mtrace_mod_mem_write_read; // @[myCPU.scala 138:29]
  wire [2:0] _mtrace_mod_mem_size; // @[myCPU.scala 138:29]
  wire  _mtrace_mod_mem_cached; // @[myCPU.scala 138:29]
  wire  fifo_with_bundle_clock; // @[myCPU.scala 159:29]
  wire  fifo_with_bundle_reset; // @[myCPU.scala 159:29]
  wire [1:0] fifo_with_bundle_io_read_en; // @[myCPU.scala 159:29]
  wire [1:0] fifo_with_bundle_io_write_en; // @[myCPU.scala 159:29]
  wire [63:0] fifo_with_bundle_io_read_out_0_pc; // @[myCPU.scala 159:29]
  wire [31:0] fifo_with_bundle_io_read_out_0_inst; // @[myCPU.scala 159:29]
  wire [1:0] fifo_with_bundle_io_read_out_0_exception_type; // @[myCPU.scala 159:29]
  wire [63:0] fifo_with_bundle_io_read_out_0_pre_pc_target; // @[myCPU.scala 159:29]
  wire [6:0] fifo_with_bundle_io_read_out_0_pre_lookup_data; // @[myCPU.scala 159:29]
  wire [3:0] fifo_with_bundle_io_read_out_0_pre_hashcode; // @[myCPU.scala 159:29]
  wire [1:0] fifo_with_bundle_io_read_out_0_pre_pht; // @[myCPU.scala 159:29]
  wire [6:0] fifo_with_bundle_io_read_out_0_pre_bht; // @[myCPU.scala 159:29]
  wire [7:0] fifo_with_bundle_io_read_out_0_pre_lookup_value; // @[myCPU.scala 159:29]
  wire  fifo_with_bundle_io_read_out_0_pre_decoder_branchD_flag; // @[myCPU.scala 159:29]
  wire  fifo_with_bundle_io_read_out_0_pre_decoder_jump; // @[myCPU.scala 159:29]
  wire [5:0] fifo_with_bundle_io_read_out_0_pre_decoder_branchdata; // @[myCPU.scala 159:29]
  wire  fifo_with_bundle_io_read_out_0_pre_decoder_jr; // @[myCPU.scala 159:29]
  wire  fifo_with_bundle_io_read_out_0_true_branch_state; // @[myCPU.scala 159:29]
  wire [63:0] fifo_with_bundle_io_write_in_0_pc; // @[myCPU.scala 159:29]
  wire [31:0] fifo_with_bundle_io_write_in_0_inst; // @[myCPU.scala 159:29]
  wire [63:0] fifo_with_bundle_io_write_in_0_pre_pc_target; // @[myCPU.scala 159:29]
  wire [6:0] fifo_with_bundle_io_write_in_0_pre_lookup_data; // @[myCPU.scala 159:29]
  wire [3:0] fifo_with_bundle_io_write_in_0_pre_hashcode; // @[myCPU.scala 159:29]
  wire [1:0] fifo_with_bundle_io_write_in_0_pre_pht; // @[myCPU.scala 159:29]
  wire [6:0] fifo_with_bundle_io_write_in_0_pre_bht; // @[myCPU.scala 159:29]
  wire [7:0] fifo_with_bundle_io_write_in_0_pre_lookup_value; // @[myCPU.scala 159:29]
  wire  fifo_with_bundle_io_write_in_0_pre_decoder_branchD_flag; // @[myCPU.scala 159:29]
  wire  fifo_with_bundle_io_write_in_0_pre_decoder_jump; // @[myCPU.scala 159:29]
  wire [5:0] fifo_with_bundle_io_write_in_0_pre_decoder_branchdata; // @[myCPU.scala 159:29]
  wire  fifo_with_bundle_io_write_in_0_pre_decoder_jr; // @[myCPU.scala 159:29]
  wire  fifo_with_bundle_io_write_in_0_true_branch_state; // @[myCPU.scala 159:29]
  wire  fifo_with_bundle_io_full; // @[myCPU.scala 159:29]
  wire  fifo_with_bundle_io_empty; // @[myCPU.scala 159:29]
  wire  fifo_with_bundle_io_point_write_en; // @[myCPU.scala 159:29]
  wire  fifo_with_bundle_io_point_flush; // @[myCPU.scala 159:29]
  wire  stage_fec_1_pc_L_clock; // @[myCPU.scala 421:34]
  wire  stage_fec_1_pc_L_reset; // @[myCPU.scala 421:34]
  wire  stage_fec_1_pc_L_io_stall; // @[myCPU.scala 421:34]
  wire  stage_fec_1_pc_L_io_flush; // @[myCPU.scala 421:34]
  wire [63:0] stage_fec_1_pc_L_io_in_pc_value_in; // @[myCPU.scala 421:34]
  wire [63:0] stage_fec_1_pc_L_io_out_pc_value_out; // @[myCPU.scala 421:34]
  wire  stage_fec_1_pc_M_clock; // @[myCPU.scala 422:34]
  wire  stage_fec_1_pc_M_reset; // @[myCPU.scala 422:34]
  wire  stage_fec_1_pc_M_io_stall; // @[myCPU.scala 422:34]
  wire  stage_fec_1_pc_M_io_flush; // @[myCPU.scala 422:34]
  wire [63:0] stage_fec_1_pc_M_io_in_pc_value_in; // @[myCPU.scala 422:34]
  wire [63:0] stage_fec_1_pc_M_io_out_pc_value_out; // @[myCPU.scala 422:34]
  wire  stage_fec_1_pc_R_clock; // @[myCPU.scala 423:34]
  wire  stage_fec_1_pc_R_reset; // @[myCPU.scala 423:34]
  wire  stage_fec_1_pc_R_io_stall; // @[myCPU.scala 423:34]
  wire  stage_fec_1_pc_R_io_flush; // @[myCPU.scala 423:34]
  wire [63:0] stage_fec_1_pc_R_io_in_pc_value_in; // @[myCPU.scala 423:34]
  wire [63:0] stage_fec_1_pc_R_io_out_pc_value_out; // @[myCPU.scala 423:34]
  wire  branch_prediction_with_blockram_clock; // @[myCPU.scala 452:21]
  wire  branch_prediction_with_blockram_reset; // @[myCPU.scala 452:21]
  wire [63:0] branch_prediction_with_blockram_io_pc; // @[myCPU.scala 452:21]
  wire [63:0] branch_prediction_with_blockram_io_write_pc; // @[myCPU.scala 452:21]
  wire [3:0] branch_prediction_with_blockram_io_aw_pht_ways_addr; // @[myCPU.scala 452:21]
  wire [6:0] branch_prediction_with_blockram_io_aw_pht_addr; // @[myCPU.scala 452:21]
  wire [6:0] branch_prediction_with_blockram_io_aw_bht_addr; // @[myCPU.scala 452:21]
  wire [63:0] branch_prediction_with_blockram_io_aw_target_addr; // @[myCPU.scala 452:21]
  wire  branch_prediction_with_blockram_io_btb_write; // @[myCPU.scala 452:21]
  wire  branch_prediction_with_blockram_io_bht_write; // @[myCPU.scala 452:21]
  wire  branch_prediction_with_blockram_io_pht_write; // @[myCPU.scala 452:21]
  wire [6:0] branch_prediction_with_blockram_io_bht_in; // @[myCPU.scala 452:21]
  wire [7:0] branch_prediction_with_blockram_io_pht_in; // @[myCPU.scala 452:21]
  wire [1:0] branch_prediction_with_blockram_io_out_L; // @[myCPU.scala 452:21]
  wire  branch_prediction_with_blockram_io_pre_L; // @[myCPU.scala 452:21]
  wire [6:0] branch_prediction_with_blockram_io_bht_L; // @[myCPU.scala 452:21]
  wire  branch_prediction_with_blockram_io_btb_hit_0; // @[myCPU.scala 452:21]
  wire [63:0] branch_prediction_with_blockram_io_pre_target_L; // @[myCPU.scala 452:21]
  wire  branch_prediction_with_blockram_io_stage2_stall; // @[myCPU.scala 452:21]
  wire  branch_prediction_with_blockram_io_stage2_flush; // @[myCPU.scala 452:21]
  wire [7:0] branch_prediction_with_blockram_io_pht_lookup_value_out; // @[myCPU.scala 452:21]
  wire [6:0] branch_prediction_with_blockram_io_lookup_data_0; // @[myCPU.scala 452:21]
  wire  stage_fec_2_pc_L_clock; // @[myCPU.scala 521:34]
  wire  stage_fec_2_pc_L_reset; // @[myCPU.scala 521:34]
  wire  stage_fec_2_pc_L_io_stall; // @[myCPU.scala 521:34]
  wire  stage_fec_2_pc_L_io_flush; // @[myCPU.scala 521:34]
  wire [63:0] stage_fec_2_pc_L_io_in_pc_value_in; // @[myCPU.scala 521:34]
  wire [63:0] stage_fec_2_pc_L_io_out_pc_value_out; // @[myCPU.scala 521:34]
  wire  stage_fec_2_pc_M_clock; // @[myCPU.scala 522:34]
  wire  stage_fec_2_pc_M_reset; // @[myCPU.scala 522:34]
  wire  stage_fec_2_pc_M_io_stall; // @[myCPU.scala 522:34]
  wire  stage_fec_2_pc_M_io_flush; // @[myCPU.scala 522:34]
  wire [63:0] stage_fec_2_pc_M_io_in_pc_value_in; // @[myCPU.scala 522:34]
  wire [63:0] stage_fec_2_pc_M_io_out_pc_value_out; // @[myCPU.scala 522:34]
  wire  stage_fec_2_pc_R_clock; // @[myCPU.scala 523:34]
  wire  stage_fec_2_pc_R_reset; // @[myCPU.scala 523:34]
  wire  stage_fec_2_pc_R_io_stall; // @[myCPU.scala 523:34]
  wire  stage_fec_2_pc_R_io_flush; // @[myCPU.scala 523:34]
  wire [63:0] stage_fec_2_pc_R_io_in_pc_value_in; // @[myCPU.scala 523:34]
  wire [63:0] stage_fec_2_pc_R_io_out_pc_value_out; // @[myCPU.scala 523:34]
  wire  id_bru_state_clock; // @[myCPU.scala 685:31]
  wire  id_bru_state_reset; // @[myCPU.scala 685:31]
  wire  id_bru_state_io_stall; // @[myCPU.scala 685:31]
  wire  id_bru_state_io_flush; // @[myCPU.scala 685:31]
  wire [1:0] id_bru_state_io_in_pht; // @[myCPU.scala 685:31]
  wire [6:0] id_bru_state_io_in_bht; // @[myCPU.scala 685:31]
  wire [3:0] id_bru_state_io_in_hashcode; // @[myCPU.scala 685:31]
  wire [63:0] id_bru_state_io_in_target_pc; // @[myCPU.scala 685:31]
  wire [6:0] id_bru_state_io_in_lookup_data; // @[myCPU.scala 685:31]
  wire [7:0] id_bru_state_io_in_pht_lookup_value; // @[myCPU.scala 685:31]
  wire [1:0] id_bru_state_io_out_pht; // @[myCPU.scala 685:31]
  wire [6:0] id_bru_state_io_out_bht; // @[myCPU.scala 685:31]
  wire [3:0] id_bru_state_io_out_hashcode; // @[myCPU.scala 685:31]
  wire [63:0] id_bru_state_io_out_target_pc; // @[myCPU.scala 685:31]
  wire [6:0] id_bru_state_io_out_lookup_data; // @[myCPU.scala 685:31]
  wire [7:0] id_bru_state_io_out_pht_lookup_value; // @[myCPU.scala 685:31]
  wire  ex_bru_state_clock; // @[myCPU.scala 689:31]
  wire  ex_bru_state_reset; // @[myCPU.scala 689:31]
  wire  ex_bru_state_io_stall; // @[myCPU.scala 689:31]
  wire  ex_bru_state_io_flush; // @[myCPU.scala 689:31]
  wire [1:0] ex_bru_state_io_in_pht; // @[myCPU.scala 689:31]
  wire [6:0] ex_bru_state_io_in_bht; // @[myCPU.scala 689:31]
  wire [3:0] ex_bru_state_io_in_hashcode; // @[myCPU.scala 689:31]
  wire [63:0] ex_bru_state_io_in_target_pc; // @[myCPU.scala 689:31]
  wire [6:0] ex_bru_state_io_in_lookup_data; // @[myCPU.scala 689:31]
  wire [7:0] ex_bru_state_io_in_pht_lookup_value; // @[myCPU.scala 689:31]
  wire [1:0] ex_bru_state_io_out_pht; // @[myCPU.scala 689:31]
  wire [6:0] ex_bru_state_io_out_bht; // @[myCPU.scala 689:31]
  wire [3:0] ex_bru_state_io_out_hashcode; // @[myCPU.scala 689:31]
  wire [63:0] ex_bru_state_io_out_target_pc; // @[myCPU.scala 689:31]
  wire [6:0] ex_bru_state_io_out_lookup_data; // @[myCPU.scala 689:31]
  wire [7:0] ex_bru_state_io_out_pht_lookup_value; // @[myCPU.scala 689:31]
  wire  mem_bru_state_clock; // @[myCPU.scala 693:32]
  wire  mem_bru_state_reset; // @[myCPU.scala 693:32]
  wire  mem_bru_state_io_stall; // @[myCPU.scala 693:32]
  wire  mem_bru_state_io_flush; // @[myCPU.scala 693:32]
  wire [1:0] mem_bru_state_io_in_pht; // @[myCPU.scala 693:32]
  wire [6:0] mem_bru_state_io_in_bht; // @[myCPU.scala 693:32]
  wire [3:0] mem_bru_state_io_in_hashcode; // @[myCPU.scala 693:32]
  wire [63:0] mem_bru_state_io_in_target_pc; // @[myCPU.scala 693:32]
  wire [6:0] mem_bru_state_io_in_lookup_data; // @[myCPU.scala 693:32]
  wire [7:0] mem_bru_state_io_in_pht_lookup_value; // @[myCPU.scala 693:32]
  wire [1:0] mem_bru_state_io_out_pht; // @[myCPU.scala 693:32]
  wire [6:0] mem_bru_state_io_out_bht; // @[myCPU.scala 693:32]
  wire [3:0] mem_bru_state_io_out_hashcode; // @[myCPU.scala 693:32]
  wire [63:0] mem_bru_state_io_out_target_pc; // @[myCPU.scala 693:32]
  wire [6:0] mem_bru_state_io_out_lookup_data; // @[myCPU.scala 693:32]
  wire [7:0] mem_bru_state_io_out_pht_lookup_value; // @[myCPU.scala 693:32]
  wire  mem2_bru_state_clock; // @[myCPU.scala 697:33]
  wire  mem2_bru_state_reset; // @[myCPU.scala 697:33]
  wire  mem2_bru_state_io_stall; // @[myCPU.scala 697:33]
  wire  mem2_bru_state_io_flush; // @[myCPU.scala 697:33]
  wire [1:0] mem2_bru_state_io_in_pht; // @[myCPU.scala 697:33]
  wire [6:0] mem2_bru_state_io_in_bht; // @[myCPU.scala 697:33]
  wire [3:0] mem2_bru_state_io_in_hashcode; // @[myCPU.scala 697:33]
  wire [63:0] mem2_bru_state_io_in_target_pc; // @[myCPU.scala 697:33]
  wire [6:0] mem2_bru_state_io_in_lookup_data; // @[myCPU.scala 697:33]
  wire [7:0] mem2_bru_state_io_in_pht_lookup_value; // @[myCPU.scala 697:33]
  wire [1:0] mem2_bru_state_io_out_pht; // @[myCPU.scala 697:33]
  wire [6:0] mem2_bru_state_io_out_bht; // @[myCPU.scala 697:33]
  wire [3:0] mem2_bru_state_io_out_hashcode; // @[myCPU.scala 697:33]
  wire [63:0] mem2_bru_state_io_out_target_pc; // @[myCPU.scala 697:33]
  wire [6:0] mem2_bru_state_io_out_lookup_data; // @[myCPU.scala 697:33]
  wire [7:0] mem2_bru_state_io_out_pht_lookup_value; // @[myCPU.scala 697:33]
  wire  wb_bru_state_clock; // @[myCPU.scala 701:31]
  wire  wb_bru_state_reset; // @[myCPU.scala 701:31]
  wire  wb_bru_state_io_stall; // @[myCPU.scala 701:31]
  wire  wb_bru_state_io_flush; // @[myCPU.scala 701:31]
  wire [1:0] wb_bru_state_io_in_pht; // @[myCPU.scala 701:31]
  wire [6:0] wb_bru_state_io_in_bht; // @[myCPU.scala 701:31]
  wire [3:0] wb_bru_state_io_in_hashcode; // @[myCPU.scala 701:31]
  wire [63:0] wb_bru_state_io_in_target_pc; // @[myCPU.scala 701:31]
  wire [6:0] wb_bru_state_io_in_lookup_data; // @[myCPU.scala 701:31]
  wire [7:0] wb_bru_state_io_in_pht_lookup_value; // @[myCPU.scala 701:31]
  wire [1:0] wb_bru_state_io_out_pht; // @[myCPU.scala 701:31]
  wire [6:0] wb_bru_state_io_out_bht; // @[myCPU.scala 701:31]
  wire [3:0] wb_bru_state_io_out_hashcode; // @[myCPU.scala 701:31]
  wire [63:0] wb_bru_state_io_out_target_pc; // @[myCPU.scala 701:31]
  wire [6:0] wb_bru_state_io_out_lookup_data; // @[myCPU.scala 701:31]
  wire [7:0] wb_bru_state_io_out_pht_lookup_value; // @[myCPU.scala 701:31]
  wire  _commit_difftest_reset; // @[myCPU.scala 1148:34]
  wire  _commit_difftest_clock; // @[myCPU.scala 1148:34]
  wire [2047:0] _commit_difftest_gpr_wire; // @[myCPU.scala 1148:34]
  wire [63:0] _commit_difftest_pc; // @[myCPU.scala 1148:34]
  wire [63:0] _commit_difftest_debug_pc; // @[myCPU.scala 1148:34]
  wire  _commit_difftest_inst_commit; // @[myCPU.scala 1148:34]
  wire  _commit_difftest_data_ok_ok; // @[myCPU.scala 1148:34]
  wire  _commit_difftest_cpu_ebreak_sign; // @[myCPU.scala 1148:34]
  wire  _T_2 = ~resetn; // @[myCPU.scala 114:41]
  wire  stage_fec_2_inst_jump = inst_sram_rdata_L[33]; // @[myCPU.scala 179:45]
  wire  stage_fec_2_inst_branch = inst_sram_rdata_L[32]; // @[myCPU.scala 180:47]
  reg  pre_decoder_branchD_flag; // @[myCPU.scala 182:44]
  reg [5:0] pre_decoder_branchdata; // @[myCPU.scala 183:43]
  reg  pre_decoder_jump; // @[myCPU.scala 184:40]
  reg  pre_decoder_jr; // @[myCPU.scala 185:40]
  wire [12:0] _immSB_T_4 = {_if2id_io_InstrD[31],_if2id_io_InstrD[7],_if2id_io_InstrD[30:25],_if2id_io_InstrD[11:8],1'h0
    }; // @[Cat.scala 31:58]
  wire [5:0] immSB_lo_lo_lo = {_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12]
    }; // @[Cat.scala 31:58]
  wire [11:0] immSB_lo_lo = {_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],
    immSB_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [12:0] immSB_lo_hi = {_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],
    _immSB_T_4[12],immSB_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [24:0] immSB_lo_1 = {_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],
    _immSB_T_4[12],immSB_lo_lo_lo,immSB_lo_lo}; // @[Cat.scala 31:58]
  wire [50:0] _immSB_T_56 = {_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],_immSB_T_4[12],
    _immSB_T_4[12],immSB_lo_lo_lo,immSB_lo_hi,immSB_lo_1}; // @[Cat.scala 31:58]
  wire [63:0] immSB = {_immSB_T_56,_if2id_io_InstrD[31],_if2id_io_InstrD[7],_if2id_io_InstrD[30:25],_if2id_io_InstrD[11:
    8],1'h0}; // @[Cat.scala 31:58]
  wire  _PCSrcD_T_1 = _cfu_io_StallD; // @[myCPU.scala 200:66]
  wire  _PCSrcD_T_3 = _br_io_exe; // @[myCPU.scala 200:85]
  wire [63:0] PCBranchD = immSB + _if2id_io_PCD; // @[myCPU.scala 201:27]
  wire [20:0] _immUJ_T_4 = {_if2id_io_InstrD[31],_if2id_io_InstrD[19:12],_if2id_io_InstrD[20],_if2id_io_InstrD[30:21],1'h0
    }; // @[Cat.scala 31:58]
  wire [4:0] immUJ_lo_lo_lo = {_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20]}; // @[Cat.scala 31:58]
  wire [9:0] immUJ_lo_lo = {_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],
    _immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20]}; // @[Cat.scala 31:58]
  wire [10:0] immUJ_lo_hi = {_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],
    immUJ_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [20:0] immUJ_lo_1 = {_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],
    immUJ_lo_lo_lo,immUJ_lo_lo}; // @[Cat.scala 31:58]
  wire [63:0] immUJ = {_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],_immUJ_T_4[20],
    immUJ_lo_lo_lo,immUJ_lo_hi,immUJ_lo_1,_immUJ_T_4}; // @[Cat.scala 31:58]
  wire [5:0] PCJumpD_lo_lo_lo = {_if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],
    _if2id_io_InstrD[31],_if2id_io_InstrD[31]}; // @[Cat.scala 31:58]
  wire [12:0] PCJumpD_lo_lo = {_if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],
    _if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],PCJumpD_lo_lo_lo}; // @[Cat.scala 31:58]
  wire [25:0] PCJumpD_lo = {_if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],
    _if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],PCJumpD_lo_lo_lo,PCJumpD_lo_lo}; // @[Cat.scala 31:58]
  wire [51:0] _PCJumpD_T_54 = {_if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],
    _if2id_io_InstrD[31],_if2id_io_InstrD[31],_if2id_io_InstrD[31],PCJumpD_lo_lo_lo,PCJumpD_lo_lo,PCJumpD_lo}; // @[Cat.scala 31:58]
  wire [63:0] _PCJumpD_T_56 = {_PCJumpD_T_54,_if2id_io_InstrD[31:20]}; // @[Cat.scala 31:58]
  reg [63:0] resultE2M_Reg; // @[myCPU.scala 981:32]
  reg [63:0] ResultM2_Reg; // @[myCPU.scala 1035:29]
  wire [63:0] _BranchR1D_T_2 = _cfu_io_Forward1D[1] ? ResultM2_Reg : _regfile_io_RD1; // @[myCPU.scala 773:61]
  wire [63:0] BranchR1D = _cfu_io_Forward1D[0] ? resultE2M_Reg : _BranchR1D_T_2; // @[myCPU.scala 773:20]
  wire [63:0] _PCJumpD_T_58 = BranchR1D + _PCJumpD_T_56; // @[myCPU.scala 204:58]
  wire [63:0] _PCJumpD_T_60 = immUJ + _if2id_io_PCD; // @[myCPU.scala 204:107]
  wire [63:0] PCJumpD = pre_decoder_jr ? _PCJumpD_T_58 : _PCJumpD_T_60; // @[myCPU.scala 204:24]
  reg [63:0] PCW_Reg; // @[myCPU.scala 292:26]
  wire  _PCW_Reg_T = _mem22wb_io_PCW != 64'h0; // @[myCPU.scala 296:36]
  reg [63:0] reg_pc; // @[myCPU.scala 301:25]
  reg  wb_exception; // @[myCPU.scala 637:31]
  wire  RegWriteW = wb_exception ? 1'h0 : _mem22wb_io_RegWriteW_Out; // @[myCPU.scala 1162:21]
  wire [3:0] _debug_wb_rf_wen_T_2 = RegWriteW ? 4'hf : 4'h0; // @[myCPU.scala 304:62]
  reg [63:0] pc_next_wait; // @[myCPU.scala 342:31]
  wire  ready_to_branch = fifo_with_bundle_io_point_write_en; // @[myCPU.scala 344:31 599:21]
  reg  stage_fec_2_stall_reg; // @[myCPU.scala 508:40]
  reg  stage_fec_2_valid; // @[myCPU.scala 479:36]
  wire  _stage_fec_2_branch_answer_T_7 = _csr_io_exception; // @[myCPU.scala 511:209]
  wire  _stage_fec_2_branch_answer_T_8 = ~_csr_io_exception; // @[myCPU.scala 511:190]
  wire  stage_fec_2_branch_answer = branch_prediction_with_blockram_io_pre_L & (stage_fec_2_inst_branch |
    stage_fec_2_inst_jump) & branch_prediction_with_blockram_io_btb_hit_0 & stage_fec_2_stall_reg & stage_fec_2_valid &
    ~_csr_io_exception; // @[myCPU.scala 511:187]
  wire  _pc_next_wait_T = ready_to_branch | stage_fec_2_branch_answer; // @[myCPU.scala 345:41]
  wire [63:0] _PC_nextD_T_2 = _PCSrcD_T_3 ? PCBranchD : _if2id_io_PCPlus4D; // @[Mux.scala 101:16]
  wire [63:0] PC_nextD = pre_decoder_jump ? PCJumpD : _PC_nextD_T_2; // @[Mux.scala 101:16]
  wire [63:0] stage_fec_2_pre_target_0 = branch_prediction_with_blockram_io_pre_target_L; // @[myCPU.scala 484:38 500:31]
  wire [63:0] stage_fec_1_pc = stage_fec_1_pc_L_io_out_pc_value_out; // @[myCPU.scala 176:26 449:20]
  wire [63:0] _stage_fec_1_pc_next_T_1 = stage_fec_1_pc + 64'h4; // @[myCPU.scala 416:93]
  wire [63:0] stage_fec_1_pc_next = stage_fec_2_branch_answer ? stage_fec_2_pre_target_0 : _stage_fec_1_pc_next_T_1; // @[myCPU.scala 416:31]
  wire [63:0] Pc_Next_normal = fifo_with_bundle_io_point_write_en ? PC_nextD : stage_fec_1_pc_next; // @[myCPU.scala 765:26]
  reg  pc_req_wait; // @[myCPU.scala 346:30]
  wire  _T_4 = ~inst_sram_en; // @[myCPU.scala 350:10]
  wire  _GEN_0 = pc_req_wait & inst_sram_en | _stage_fec_2_branch_answer_T_7 | ready_to_branch & inst_sram_en ? 1'h0 :
    pc_req_wait; // @[myCPU.scala 352:119 353:21 355:21]
  reg [63:0] exception_Pc_reg; // @[myCPU.scala 359:35]
  reg  returnPc_req_wait; // @[myCPU.scala 362:36]
  wire  _GEN_2 = returnPc_req_wait & inst_sram_en ? 1'h0 : returnPc_req_wait; // @[myCPU.scala 367:54 368:27 370:27]
  wire [63:0] _Pc_Next_T_1 = pc_req_wait ? pc_next_wait : Pc_Next_normal; // @[myCPU.scala 377:140]
  wire [63:0] _Pc_Next_T_2 = ready_to_branch ? Pc_Next_normal : _Pc_Next_T_1; // @[myCPU.scala 377:105]
  wire [63:0] _Pc_Next_T_3 = returnPc_req_wait ? exception_Pc_reg : _Pc_Next_T_2; // @[myCPU.scala 377:66]
  wire [63:0] Pc_Next = _stage_fec_2_branch_answer_T_7 ? _csr_io_return_pc : _Pc_Next_T_3; // @[myCPU.scala 377:19]
  wire  _commit_cache_reg_T = _cfu_io_StallE; // @[myCPU.scala 399:40]
  reg  stage_fec_1_valid; // @[myCPU.scala 458:36]
  wire  _stage_fec_1_valid_T_2 = _pc_next_wait_T ? 1'h0 : stage_fec_1_valid; // @[myCPU.scala 462:55]
  wire  stage_fec_2_stall = stage2_stall & ~_pc_next_wait_T; // @[myCPU.scala 472:42]
  reg [6:0] stage_fec_2_bht_0; // @[myCPU.scala 482:35]
  reg [3:0] stage_fec_2_hascode_0; // @[myCPU.scala 486:39]
  wire  stage_fec_2_hascode_0_num_array_0 = ^branch_prediction_with_blockram_io_pc[7:4]; // @[macros.scala 447:45]
  wire  stage_fec_2_hascode_0_num_array_1 = ^branch_prediction_with_blockram_io_pc[11:8]; // @[macros.scala 447:45]
  wire  stage_fec_2_hascode_0_num_array_2 = ^branch_prediction_with_blockram_io_pc[15:12]; // @[macros.scala 447:45]
  wire  stage_fec_2_hascode_0_num_array_3 = ^branch_prediction_with_blockram_io_pc[19:16]; // @[macros.scala 447:45]
  wire [3:0] _stage_fec_2_hascode_0_T_1 = {stage_fec_2_hascode_0_num_array_3,stage_fec_2_hascode_0_num_array_2,
    stage_fec_2_hascode_0_num_array_1,stage_fec_2_hascode_0_num_array_0}; // @[macros.scala 449:13]
  wire  _stage_fec_2_data_valid_T = ~fifo_with_bundle_io_empty; // @[myCPU.scala 529:88]
  wire [31:0] inst_buffer_write_bundle_inst = inst_sram_rdata_L[31:0]; // @[myCPU.scala 551:60]
  wire [6:0] inst_buffer_write_bundle_pre_decoder_jr_opD = inst_buffer_write_bundle_inst[6:0]; // @[macros.scala 495:24]
  wire [2:0] inst_buffer_write_bundle_pre_decoder_jr_Funct3D = inst_buffer_write_bundle_inst[14:12]; // @[macros.scala 496:28]
  wire  _T_25 = _cfu_io_StallF; // @[myCPU.scala 577:51]
  wire  _pre_decoder_branchD_flag_T = _cfu_io_FlushD; // @[myCPU.scala 606:52]
  wire  inst_buffer_read_out_pre_decoder_branchD_flag = fifo_with_bundle_io_read_out_0_pre_decoder_branchD_flag; // @[myCPU.scala 602:36 603:26]
  wire  inst_buffer_read_out_pre_decoder_jump = fifo_with_bundle_io_read_out_0_pre_decoder_jump; // @[myCPU.scala 602:36 603:26]
  wire [5:0] inst_buffer_read_out_pre_decoder_branchdata = fifo_with_bundle_io_read_out_0_pre_decoder_branchdata; // @[myCPU.scala 602:36 603:26]
  wire  inst_buffer_read_out_pre_decoder_jr = fifo_with_bundle_io_read_out_0_pre_decoder_jr; // @[myCPU.scala 602:36 603:26]
  wire  __if2id_io_InstrF_T = _cu_io1_BadInstrD; // @[myCPU.scala 621:52]
  wire  __if2id_io_InstrF_T_1 = _cu_io1_SysCallD; // @[myCPU.scala 621:79]
  wire  __if2id_io_InstrF_T_3 = _cu_io1_EretD; // @[myCPU.scala 622:47]
  wire [31:0] inst_buffer_read_out_inst = fifo_with_bundle_io_read_out_0_inst; // @[myCPU.scala 602:36 603:26]
  wire [31:0] __if2id_io_InstrF_T_5 = _cu_io1_BadInstrD | _cu_io1_SysCallD | __if2id_io_InstrF_T_3 ? 32'h0 :
    inst_buffer_read_out_inst; // @[myCPU.scala 621:33]
  reg  id_exception; // @[myCPU.scala 625:31]
  wire [63:0] inst_buffer_read_out_pc = fifo_with_bundle_io_read_out_0_pc; // @[myCPU.scala 602:36 603:26]
  wire [1:0] inst_buffer_read_out_exception_type = fifo_with_bundle_io_read_out_0_exception_type; // @[myCPU.scala 602:36 603:26]
  reg  ex_exception; // @[myCPU.scala 628:31]
  wire  _ex_exception_T = _cfu_io_FlushE; // @[myCPU.scala 629:40]
  reg  mem_exception; // @[myCPU.scala 631:32]
  wire  _mem_exception_T = _cfu_io_FlushM; // @[myCPU.scala 632:41]
  wire  _mem_exception_T_1 = _cfu_io_StallM; // @[myCPU.scala 632:71]
  reg  mem2_exception; // @[myCPU.scala 634:33]
  wire  _mem2_exception_T = _cfu_io_FlushM2; // @[myCPU.scala 635:43]
  wire  _mem2_exception_T_1 = _cfu_io_StallM2; // @[myCPU.scala 635:74]
  wire  _wb_exception_T = _cfu_io_FlushW; // @[myCPU.scala 638:40]
  wire  _wb_exception_T_1 = _cfu_io_StallW; // @[myCPU.scala 638:70]
  reg  id_true_branch_state; // @[myCPU.scala 682:39]
  wire  inst_buffer_read_out_true_branch_state = fifo_with_bundle_io_read_out_0_true_branch_state; // @[myCPU.scala 602:36 603:26]
  reg  inst_tlb_exceptionE; // @[myCPU.scala 712:38]
  wire  target_neq_branchD = id_bru_state_io_out_target_pc != PCBranchD; // @[myCPU.scala 726:62]
  wire  target_neq_jumpD = id_bru_state_io_out_target_pc != PCJumpD; // @[myCPU.scala 727:62]
  wire  target_addr_error = pre_decoder_jump & target_neq_jumpD | _PCSrcD_T_3 & target_neq_branchD; // @[myCPU.scala 729:75]
  wire  _T_31 = pre_decoder_jump | _PCSrcD_T_3; // @[myCPU.scala 732:117]
  wire  _T_37 = ex_exception | mem_exception | mem2_exception | wb_exception; // @[myCPU.scala 732:241]
  wire [63:0] _Pc_targetD_T_2 = pre_decoder_jump ? PCJumpD : 64'h0; // @[Mux.scala 101:16]
  reg  true_branch_stateE; // @[myCPU.scala 743:37]
  wire [1:0] _pht_tobeE_T_1 = true_branch_stateE ? 2'h3 : 2'h2; // @[macros.scala 468:30]
  wire [1:0] _pht_tobeE_T_2 = true_branch_stateE ? 2'h2 : 2'h0; // @[macros.scala 469:32]
  wire [1:0] _pht_tobeE_T_3 = true_branch_stateE ? 2'h3 : 2'h1; // @[macros.scala 470:30]
  wire [1:0] _pht_tobeE_T_5 = 2'h3 == ex_bru_state_io_out_pht ? _pht_tobeE_T_1 : {{1'd0}, true_branch_stateE}; // @[Mux.scala 81:58]
  wire [1:0] _pht_tobeE_T_7 = 2'h1 == ex_bru_state_io_out_pht ? _pht_tobeE_T_2 : _pht_tobeE_T_5; // @[Mux.scala 81:58]
  wire [1:0] pht_tobeE = 2'h2 == ex_bru_state_io_out_pht ? _pht_tobeE_T_3 : _pht_tobeE_T_7; // @[Mux.scala 81:58]
  wire [7:0] _pht_lookup_value_tobeE_T_2 = {ex_bru_state_io_out_pht_lookup_value[7:2],pht_tobeE}; // @[Cat.scala 31:58]
  wire [7:0] _pht_lookup_value_tobeE_T_5 = {ex_bru_state_io_out_pht_lookup_value[7:4],pht_tobeE,
    ex_bru_state_io_out_pht_lookup_value[1:0]}; // @[Cat.scala 31:58]
  wire [7:0] _pht_lookup_value_tobeE_T_8 = {ex_bru_state_io_out_pht_lookup_value[7:6],pht_tobeE,
    ex_bru_state_io_out_pht_lookup_value[3:0]}; // @[Cat.scala 31:58]
  wire [7:0] _pht_lookup_value_tobeE_T_10 = {pht_tobeE,ex_bru_state_io_out_pht_lookup_value[5:0]}; // @[Cat.scala 31:58]
  wire [7:0] _pht_lookup_value_tobeE_T_12 = 2'h1 == ex_bru_state_io_out_lookup_data[1:0] ? _pht_lookup_value_tobeE_T_5
     : _pht_lookup_value_tobeE_T_2; // @[Mux.scala 81:58]
  wire [7:0] _pht_lookup_value_tobeE_T_14 = 2'h2 == ex_bru_state_io_out_lookup_data[1:0] ? _pht_lookup_value_tobeE_T_8
     : _pht_lookup_value_tobeE_T_12; // @[Mux.scala 81:58]
  wire [63:0] _BranchR2D_T_2 = _cfu_io_Forward2D[1] ? ResultM2_Reg : _regfile_io_RD2; // @[myCPU.scala 775:61]
  wire  _ExceptionTypeD_Out_T_1 = _if2id_io_PCD[1:0] != 2'h0; // @[myCPU.scala 777:29]
  wire [20:0] _ExceptionTypeD_Out_T_4 = _ExceptionTypeD_Out_T_1 ? 21'h100000 : 21'h0; // @[Mux.scala 27:73]
  wire [3:0] _ExceptionTypeD_Out_T_5 = _if2id_io_ExceptionTypeD_Out[0] ? 4'h8 : 4'h0; // @[Mux.scala 27:73]
  wire [2:0] _ExceptionTypeD_Out_T_6 = _if2id_io_ExceptionTypeD_Out[1] ? 3'h4 : 3'h0; // @[Mux.scala 27:73]
  wire [24:0] _ExceptionTypeD_Out_T_7 = _cu_io_fence_i_control ? 25'h1000000 : 25'h0; // @[Mux.scala 27:73]
  wire [20:0] _GEN_12 = {{17'd0}, _ExceptionTypeD_Out_T_5}; // @[Mux.scala 27:73]
  wire [20:0] _ExceptionTypeD_Out_T_8 = _ExceptionTypeD_Out_T_4 | _GEN_12; // @[Mux.scala 27:73]
  wire [20:0] _GEN_13 = {{18'd0}, _ExceptionTypeD_Out_T_6}; // @[Mux.scala 27:73]
  wire [20:0] _ExceptionTypeD_Out_T_9 = _ExceptionTypeD_Out_T_8 | _GEN_13; // @[Mux.scala 27:73]
  wire [24:0] _GEN_14 = {{4'd0}, _ExceptionTypeD_Out_T_9}; // @[Mux.scala 27:73]
  wire [24:0] _ExceptionTypeD_Out_T_10 = _GEN_14 | _ExceptionTypeD_Out_T_7; // @[Mux.scala 27:73]
  reg  int_instanceE_timer; // @[myCPU.scala 786:33]
  reg  int_instanceM_timer; // @[myCPU.scala 787:33]
  reg  int_instanceM2_timer; // @[myCPU.scala 788:33]
  reg  int_instanceW_timer; // @[myCPU.scala 789:33]
  wire [63:0] ExceptionTypeD_Out = {{39'd0}, _ExceptionTypeD_Out_T_10}; // @[myCPU.scala 192:34 776:24]
  wire [10:0] __id2ex_io_ExceptionTypeD_T_5 = __if2id_io_InstrF_T ? 11'h400 : 11'h0; // @[myCPU.scala 803:13]
  wire [8:0] __id2ex_io_ExceptionTypeD_T_7 = __if2id_io_InstrF_T_1 ? 9'h100 : 9'h0; // @[myCPU.scala 804:13]
  wire [10:0] _GEN_15 = {{2'd0}, __id2ex_io_ExceptionTypeD_T_7}; // @[myCPU.scala 803:59]
  wire [10:0] __id2ex_io_ExceptionTypeD_T_8 = __id2ex_io_ExceptionTypeD_T_5 | _GEN_15; // @[myCPU.scala 803:59]
  wire [31:0] __id2ex_io_ExceptionTypeD_T_10 = __if2id_io_InstrF_T_3 ? 32'h80000000 : 32'h0; // @[myCPU.scala 806:13]
  wire [31:0] _GEN_16 = {{21'd0}, __id2ex_io_ExceptionTypeD_T_8}; // @[myCPU.scala 804:59]
  wire [31:0] __id2ex_io_ExceptionTypeD_T_11 = _GEN_16 | __id2ex_io_ExceptionTypeD_T_10; // @[myCPU.scala 804:59]
  wire [63:0] __id2ex_io_ExceptionTypeD_T_12 = ExceptionTypeD_Out == 64'h0 ? {{32'd0}, __id2ex_io_ExceptionTypeD_T_11}
     : ExceptionTypeD_Out; // @[myCPU.scala 802:129]
  wire [63:0] __id2ex_io_ExceptionTypeD_T_13 = ext_int_timer & _csr_io_int_type_able_timer & _csr_io_Int_able ? 64'h1 :
    __id2ex_io_ExceptionTypeD_T_12; // @[myCPU.scala 802:37]
  wire  __id2ex_io_BranchJump_JrD_T_2 = pre_decoder_branchD_flag | pre_decoder_jump; // @[myCPU.scala 828:79]
  reg  inst_tlb_exceptionM; // @[myCPU.scala 841:34]
  wire [63:0] ResultW = _mem22wb_io_ResultW; // @[myCPU.scala 1161:15 289:26]
  wire [63:0] _RD1ForWardE_p_T_1 = 2'h1 == _cfu_io_Forward1E ? ResultW : _id2ex_io_RD1E; // @[Mux.scala 81:58]
  wire [63:0] _RD1ForWardE_p_T_3 = 2'h2 == _cfu_io_Forward1E ? resultE2M_Reg : _RD1ForWardE_p_T_1; // @[Mux.scala 81:58]
  wire [63:0] RD1ForWardE_p = 2'h3 == _cfu_io_Forward1E ? ResultM2_Reg : _RD1ForWardE_p_T_3; // @[Mux.scala 81:58]
  wire [63:0] _RD2ForWardE_p_T_1 = 2'h1 == _cfu_io_Forward2E ? ResultW : _id2ex_io_RD2E; // @[Mux.scala 81:58]
  wire [63:0] _RD2ForWardE_p_T_3 = 2'h2 == _cfu_io_Forward2E ? resultE2M_Reg : _RD2ForWardE_p_T_1; // @[Mux.scala 81:58]
  wire [63:0] RD2ForWardE_p = 2'h3 == _cfu_io_Forward2E ? ResultM2_Reg : _RD2ForWardE_p_T_3; // @[Mux.scala 81:58]
  reg [63:0] RD1ForWardE_r; // @[myCPU.scala 846:34]
  reg [63:0] RD2ForWardE_r; // @[myCPU.scala 847:34]
  reg  Forward_Lock1E; // @[myCPU.scala 848:34]
  reg  Forward_Lock2E; // @[myCPU.scala 849:34]
  wire [63:0] _Forward_csr_data_T_1 = 2'h1 == _cfu_io_ForwardcsrE ? _ex2mem_io_WriteDataM : _csr_io_csr_read_data; // @[Mux.scala 81:58]
  wire [63:0] Forward_csr_data = 2'h2 == _cfu_io_ForwardcsrE ? _mem2mem2_io_WriteDataM : _Forward_csr_data_T_1; // @[Mux.scala 81:58]
  wire [63:0] RD1ForWardE = Forward_Lock1E ? RD1ForWardE_r : RD1ForWardE_p; // @[myCPU.scala 854:23]
  wire [63:0] RD2ForWardE = Forward_Lock2E ? RD2ForWardE_r : RD2ForWardE_p; // @[myCPU.scala 855:23]
  wire  _Forward_Lock1E_T = _ex2mem_io_MemToRegM; // @[myCPU.scala 861:54]
  wire  _Forward_Lock1E_T_1 = _mem2mem2_io_MemToRegM; // @[myCPU.scala 861:87]
  wire  _Forward_Lock1E_T_3 = ~(_ex2mem_io_MemToRegM | _mem2mem2_io_MemToRegM); // @[myCPU.scala 861:31]
  wire [63:0] Src1E = _id2ex_io2_ALUSrcE_0 ? _id2ex_io2_PCE : RD1ForWardE; // @[myCPU.scala 876:20]
  wire [63:0] Src2E = _id2ex_io2_ALUSrcE_1 ? _id2ex_io_ImmE : RD2ForWardE; // @[myCPU.scala 883:20]
  wire  csrToRegE = _id2ex_io_ExceptionTypeE_Out == 32'h0 & _id2ex_io_csrToRegE_Out; // @[myCPU.scala 887:24]
  wire  __muldiv_io_en_T_2 = _ex2mem_io_RegWriteM; // @[myCPU.scala 894:105]
  wire  __muldiv_io_en_T_10 = _id2ex_io_R1E == _ex2mem_io_WriteRegM & __muldiv_io_en_T_2 & _Forward_Lock1E_T; // @[myCPU.scala 895:88]
  wire  __muldiv_io_en_T_11 = _id2ex_io_R2E == _ex2mem_io_WriteRegM & _ex2mem_io_RegWriteM & _Forward_Lock1E_T |
    __muldiv_io_en_T_10; // @[myCPU.scala 894:144]
  wire  __muldiv_io_en_T_13 = _mem2mem2_io_RegWriteM; // @[myCPU.scala 896:85]
  wire  __muldiv_io_en_T_16 = _id2ex_io_R2E == _mem2mem2_io_WriteRegM & _mem2mem2_io_RegWriteM & _Forward_Lock1E_T_1; // @[myCPU.scala 896:92]
  wire  __muldiv_io_en_T_17 = __muldiv_io_en_T_11 | __muldiv_io_en_T_16; // @[myCPU.scala 895:120]
  wire  __muldiv_io_en_T_22 = _id2ex_io_R1E == _mem2mem2_io_WriteRegM & __muldiv_io_en_T_13 & _Forward_Lock1E_T_1; // @[myCPU.scala 897:92]
  wire  __muldiv_io_en_T_23 = __muldiv_io_en_T_17 | __muldiv_io_en_T_22; // @[myCPU.scala 896:126]
  wire [12:0] _temp_exceptionE_T_11 = _alu_io_overflow ? 13'h1000 : 13'h0; // @[myCPU.scala 929:13]
  wire [4:0] _csr_src1_T = _id2ex_io_R1E; // @[macros.scala 435:38]
  wire [5:0] _csr_src1_T_1 = {1'h0,_csr_src1_T}; // @[Cat.scala 31:58]
  wire [63:0] csr_src1 = _id2ex_io_csr_ImmE ? {{58'd0}, _csr_src1_T_1} : RD1ForWardE; // @[myCPU.scala 959:20]
  wire [5:0] _CalCsrDataE_T = _id2ex_io_csr_controlE; // @[myCPU.scala 962:31]
  wire [63:0] _CalCsrDataE_T_2 = Forward_csr_data | csr_src1; // @[myCPU.scala 962:64]
  wire [5:0] _CalCsrDataE_T_3 = {{1'd0}, _id2ex_io_csr_controlE[5:1]}; // @[myCPU.scala 963:31]
  wire [63:0] _CalCsrDataE_T_5 = ~csr_src1; // @[myCPU.scala 963:68]
  wire [63:0] _CalCsrDataE_T_6 = Forward_csr_data & _CalCsrDataE_T_5; // @[myCPU.scala 963:64]
  wire [5:0] _CalCsrDataE_T_7 = {{2'd0}, _id2ex_io_csr_controlE[5:2]}; // @[myCPU.scala 964:31]
  wire [63:0] _CalCsrDataE_T_9 = _CalCsrDataE_T[0] ? _CalCsrDataE_T_2 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _CalCsrDataE_T_10 = _CalCsrDataE_T_3[0] ? _CalCsrDataE_T_6 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _CalCsrDataE_T_11 = _CalCsrDataE_T_7[0] ? csr_src1 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _CalCsrDataE_T_12 = _CalCsrDataE_T_9 | _CalCsrDataE_T_10; // @[Mux.scala 27:73]
  wire [63:0] CalCsrDataE = _CalCsrDataE_T_12 | _CalCsrDataE_T_11; // @[Mux.scala 27:73]
  wire  _resultE_T_1 = _id2ex_io2_LinkE; // @[myCPU.scala 977:25]
  wire [63:0] _resultE_T_2 = _id2ex_io_alu_calE ? _alu_io_result : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _resultE_T_3 = csrToRegE ? CalCsrDataE : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _resultE_T_4 = _resultE_T_1 ? _id2ex_io2_PCPlus4E : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _resultE_T_5 = _id2ex_io_muldiv_calE ? _muldiv_io_data_out : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _resultE_T_6 = _resultE_T_2 | _resultE_T_3; // @[Mux.scala 27:73]
  wire [63:0] _resultE_T_7 = _resultE_T_6 | _resultE_T_4; // @[Mux.scala 27:73]
  wire [63:0] resultE = _resultE_T_7 | _resultE_T_5; // @[Mux.scala 27:73]
  wire  __mem2mem2_io_csrWriteE_T = _ex2mem_io_csrWriteM; // @[myCPU.scala 1049:48]
  reg  tlb_exception_csr_writeM2; // @[myCPU.scala 1083:40]
  reg  tlb_exception_co0_writeW; // @[myCPU.scala 1084:40]
  wire [31:0] _Mem_withRL_Data_T_25 = {_mem2mem2_io_RtM[31:8],_dmem_io_RD[31:24]}; // @[Cat.scala 31:58]
  wire [31:0] _Mem_withRL_Data_T_22 = {_mem2mem2_io_RtM[31:16],_dmem_io_RD[31:16]}; // @[Cat.scala 31:58]
  wire [31:0] _Mem_withRL_Data_T_19 = {_mem2mem2_io_RtM[31:24],_dmem_io_RD[31:8]}; // @[Cat.scala 31:58]
  wire [63:0] _Mem_withRL_Data_T_27 = 2'h1 == _mem2mem2_io_PhyAddrM[1:0] ? {{32'd0}, _Mem_withRL_Data_T_19} :
    _dmem_io_RD; // @[Mux.scala 81:58]
  wire [63:0] _Mem_withRL_Data_T_29 = 2'h2 == _mem2mem2_io_PhyAddrM[1:0] ? {{32'd0}, _Mem_withRL_Data_T_22} :
    _Mem_withRL_Data_T_27; // @[Mux.scala 81:58]
  wire [63:0] _Mem_withRL_Data_T_31 = 2'h3 == _mem2mem2_io_PhyAddrM[1:0] ? {{32'd0}, _Mem_withRL_Data_T_25} :
    _Mem_withRL_Data_T_29; // @[Mux.scala 81:58]
  wire [31:0] _Mem_withRL_Data_T_9 = {_dmem_io_RD[23:0],_mem2mem2_io_RtM[7:0]}; // @[Cat.scala 31:58]
  wire [31:0] _Mem_withRL_Data_T_6 = {_dmem_io_RD[15:0],_mem2mem2_io_RtM[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _Mem_withRL_Data_T_3 = {_dmem_io_RD[7:0],_mem2mem2_io_RtM[23:0]}; // @[Cat.scala 31:58]
  wire [63:0] _Mem_withRL_Data_T_11 = 2'h0 == _mem2mem2_io_PhyAddrM[1:0] ? {{32'd0}, _Mem_withRL_Data_T_3} : _dmem_io_RD
    ; // @[Mux.scala 81:58]
  wire [63:0] _Mem_withRL_Data_T_13 = 2'h1 == _mem2mem2_io_PhyAddrM[1:0] ? {{32'd0}, _Mem_withRL_Data_T_6} :
    _Mem_withRL_Data_T_11; // @[Mux.scala 81:58]
  wire [63:0] _Mem_withRL_Data_T_15 = 2'h2 == _mem2mem2_io_PhyAddrM[1:0] ? {{32'd0}, _Mem_withRL_Data_T_9} :
    _Mem_withRL_Data_T_13; // @[Mux.scala 81:58]
  wire [63:0] _Mem_withRL_Data_T_33 = 2'h2 == _mem2mem2_io_MemRLM ? _Mem_withRL_Data_T_15 : _dmem_io_RD; // @[Mux.scala 81:58]
  wire [63:0] Mem_withRL_Data = 2'h1 == _mem2mem2_io_MemRLM ? _Mem_withRL_Data_T_31 : _Mem_withRL_Data_T_33; // @[Mux.scala 81:58]
  wire [63:0] __mem22wb_io_Mem_trace_budleM_data_T_2 = _mem2mem2_io_mem_trace_budleM_mem_fetch_type[0] ?
    _mem2mem2_io_mem_trace_budleM_data : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] __mem22wb_io_Mem_trace_budleM_data_T_3 = _mem2mem2_io_mem_trace_budleM_mem_fetch_type[1] ? Mem_withRL_Data
     : 64'h0; // @[Mux.scala 27:73]
  reg [63:0] pcw_reg; // @[myCPU.scala 1146:26]
  wire  csrWriteW = wb_exception ? 1'h0 : _mem22wb_io_csrWriteW; // @[myCPU.scala 1164:25]
  alu _alu ( // @[myCPU.scala 120:22]
    .io_ctrl(_alu_io_ctrl),
    .io_in1(_alu_io_in1),
    .io_in2(_alu_io_in2),
    .io_result(_alu_io_result),
    .io_overflow(_alu_io_overflow),
    .io_data_w(_alu_io_data_w)
  );
  br _br ( // @[myCPU.scala 121:22]
    .reset(_br_reset),
    .io_r1(_br_io_r1),
    .io_r2(_br_io_r2),
    .io_branch(_br_io_branch),
    .io_exe(_br_io_exe)
  );
  cfu _cfu ( // @[myCPU.scala 122:22]
    .reset(_cfu_reset),
    .io_Inst_Fifo_Empty(_cfu_io_Inst_Fifo_Empty),
    .io_dmem_calD(_cfu_io_dmem_calD),
    .io_BranchD_Flag(_cfu_io_BranchD_Flag),
    .io_JRD(_cfu_io_JRD),
    .io_CanBranchD(_cfu_io_CanBranchD),
    .io_DivPendingE(_cfu_io_DivPendingE),
    .io_DataPendingM(_cfu_io_DataPendingM),
    .io_InException(_cfu_io_InException),
    .io_WriteRegE(_cfu_io_WriteRegE),
    .io_RegWriteE(_cfu_io_RegWriteE),
    .io_csrToRegE(_cfu_io_csrToRegE),
    .io_WriteRegM(_cfu_io_WriteRegM),
    .io_MemToRegM(_cfu_io_MemToRegM),
    .io_RegWriteM(_cfu_io_RegWriteM),
    .io_csrWriteM(_cfu_io_csrWriteM),
    .io_WriteRegM2(_cfu_io_WriteRegM2),
    .io_MemToRegM2(_cfu_io_MemToRegM2),
    .io_RegWriteM2(_cfu_io_RegWriteM2),
    .io_csrWriteM2(_cfu_io_csrWriteM2),
    .io_WriteRegW(_cfu_io_WriteRegW),
    .io_RegWriteW(_cfu_io_RegWriteW),
    .io_ReadcsrAddrE(_cfu_io_ReadcsrAddrE),
    .io_WritecsrAddrM(_cfu_io_WritecsrAddrM),
    .io_WritecsrAddrM2(_cfu_io_WritecsrAddrM2),
    .io_R2D(_cfu_io_R2D),
    .io_R1D(_cfu_io_R1D),
    .io_R2E(_cfu_io_R2E),
    .io_R1E(_cfu_io_R1E),
    .io_StallF(_cfu_io_StallF),
    .io_StallD(_cfu_io_StallD),
    .io_StallE(_cfu_io_StallE),
    .io_StallM(_cfu_io_StallM),
    .io_StallM2(_cfu_io_StallM2),
    .io_StallW(_cfu_io_StallW),
    .io_FlushD(_cfu_io_FlushD),
    .io_FlushE(_cfu_io_FlushE),
    .io_FlushM(_cfu_io_FlushM),
    .io_FlushM2(_cfu_io_FlushM2),
    .io_FlushW(_cfu_io_FlushW),
    .io_Forward1E(_cfu_io_Forward1E),
    .io_Forward2E(_cfu_io_Forward2E),
    .io_Forward1D(_cfu_io_Forward1D),
    .io_Forward2D(_cfu_io_Forward2D),
    .io_ForwardcsrE(_cfu_io_ForwardcsrE)
  );
  csr _csr ( // @[myCPU.scala 123:22]
    .clock(_csr_clock),
    .reset(_csr_reset),
    .io_csr_read_addr(_csr_io_csr_read_addr),
    .io_csr_write_addr(_csr_io_csr_write_addr),
    .io_csr_write_data(_csr_io_csr_write_data),
    .io_csr_write_en(_csr_io_csr_write_en),
    .io_pc(_csr_io_pc),
    .io_exception_type_i(_csr_io_exception_type_i),
    .io_return_pc(_csr_io_return_pc),
    .io_exception(_csr_io_exception),
    .io_csr_read_data(_csr_io_csr_read_data),
    .io_icache_tags_flush(_csr_io_icache_tags_flush),
    .io_int_type_timer(_csr_io_int_type_timer),
    .io_Int_able(_csr_io_Int_able),
    .io_int_type_able_timer(_csr_io_int_type_able_timer)
  );
  cu _cu ( // @[myCPU.scala 124:22]
    .io1_InstrD(_cu_io1_InstrD),
    .io1_BadInstrD(_cu_io1_BadInstrD),
    .io1_SysCallD(_cu_io1_SysCallD),
    .io1_EretD(_cu_io1_EretD),
    .io1_dmem_addr_cal(_cu_io1_dmem_addr_cal),
    .io_RegWriteD(_cu_io_RegWriteD),
    .io_MemToRegD(_cu_io_MemToRegD),
    .io_MemWriteD(_cu_io_MemWriteD),
    .io_ALUCtrlD(_cu_io_ALUCtrlD),
    .io_ALUSrcD_0(_cu_io_ALUSrcD_0),
    .io_ALUSrcD_1(_cu_io_ALUSrcD_1),
    .io_RegDstD(_cu_io_RegDstD),
    .io_LinkD(_cu_io_LinkD),
    .io_csrWriteD(_cu_io_csrWriteD),
    .io_csrToRegD(_cu_io_csrToRegD),
    .io_LoadUnsignedD(_cu_io_LoadUnsignedD),
    .io_MemWidthD(_cu_io_MemWidthD),
    .io_ImmD(_cu_io_ImmD),
    .io_ebreakD(_cu_io_ebreakD),
    .io_data_wD(_cu_io_data_wD),
    .io_muldiv_control(_cu_io_muldiv_control),
    .io_muldiv_cal(_cu_io_muldiv_cal),
    .io_alu_cal(_cu_io_alu_cal),
    .io_csr_control(_cu_io_csr_control),
    .io_csr_Imm(_cu_io_csr_Imm),
    .io_fence_i_control(_cu_io_fence_i_control)
  );
  dmem _dmem ( // @[myCPU.scala 125:23]
    .io_data_ok(_dmem_io_data_ok),
    .io_rdata(_dmem_io_rdata),
    .io_Physisc_Address(_dmem_io_Physisc_Address),
    .io_WIDTH(_dmem_io_WIDTH),
    .io_SIGN(_dmem_io_SIGN),
    .io_RD(_dmem_io_RD),
    .io_data_pending(_dmem_io_data_pending)
  );
  dmemreq _dmemreq ( // @[myCPU.scala 126:26]
    .io_en(_dmemreq_io_en),
    .io_MemWriteE(_dmemreq_io_MemWriteE),
    .io_MemToRegE(_dmemreq_io_MemToRegE),
    .io_MemWidthE(_dmemreq_io_MemWidthE),
    .io_VAddrE(_dmemreq_io_VAddrE),
    .io_WriteDataE(_dmemreq_io_WriteDataE),
    .io_req(_dmemreq_io_req),
    .io_wr(_dmemreq_io_wr),
    .io_size(_dmemreq_io_size),
    .io_addr(_dmemreq_io_addr),
    .io_wdata(_dmemreq_io_wdata),
    .io_wstrb(_dmemreq_io_wstrb)
  );
  ex2mem _ex2mem ( // @[myCPU.scala 127:26]
    .clock(_ex2mem_clock),
    .reset(_ex2mem_reset),
    .io1_RegWriteE(_ex2mem_io1_RegWriteE),
    .io1_MemToRegE(_ex2mem_io1_MemToRegE),
    .io1_LoadUnsignedE(_ex2mem_io1_LoadUnsignedE),
    .io1_MemWidthE(_ex2mem_io1_MemWidthE),
    .io1_csrWriteE(_ex2mem_io1_csrWriteE),
    .io1_WritecsrAddrE(_ex2mem_io1_WritecsrAddrE),
    .io1_PCE(_ex2mem_io1_PCE),
    .io1_MemRLE(_ex2mem_io1_MemRLE),
    .io1_BranchJump_JrE(_ex2mem_io1_BranchJump_JrE),
    .io1_Tlb_Control(_ex2mem_io1_Tlb_Control),
    .io1_eBreakE(_ex2mem_io1_eBreakE),
    .io1_fence_i_control(_ex2mem_io1_fence_i_control),
    .io_en(_ex2mem_io_en),
    .io_clr(_ex2mem_io_clr),
    .io_WriteDataE(_ex2mem_io_WriteDataE),
    .io_WriteRegE(_ex2mem_io_WriteRegE),
    .io_PhyAddrE(_ex2mem_io_PhyAddrE),
    .io_CsrWritedataE(_ex2mem_io_CsrWritedataE),
    .io_ExceptionTypeE(_ex2mem_io_ExceptionTypeE),
    .io_RtE(_ex2mem_io_RtE),
    .io_Pc_NextE(_ex2mem_io_Pc_NextE),
    .io_mem_trace_budleE_pc(_ex2mem_io_mem_trace_budleE_pc),
    .io_mem_trace_budleE_data(_ex2mem_io_mem_trace_budleE_data),
    .io_mem_trace_budleE_mem_fetch_type(_ex2mem_io_mem_trace_budleE_mem_fetch_type),
    .io_mem_trace_budleE_addr(_ex2mem_io_mem_trace_budleE_addr),
    .io_mem_trace_budleE_len(_ex2mem_io_mem_trace_budleE_len),
    .io_mem_trace_budleE_cache(_ex2mem_io_mem_trace_budleE_cache),
    .io_RegWriteM(_ex2mem_io_RegWriteM),
    .io_MemToRegM(_ex2mem_io_MemToRegM),
    .io_WriteDataM(_ex2mem_io_WriteDataM),
    .io_WriteRegM(_ex2mem_io_WriteRegM),
    .io_LoadUnsignedM(_ex2mem_io_LoadUnsignedM),
    .io_MemWidthM(_ex2mem_io_MemWidthM),
    .io_PhyAddrM(_ex2mem_io_PhyAddrM),
    .io_csrWriteM(_ex2mem_io_csrWriteM),
    .io_WritecsrAddrM(_ex2mem_io_WritecsrAddrM),
    .io_PCM(_ex2mem_io_PCM),
    .io_ExceptionTypeM_Out(_ex2mem_io_ExceptionTypeM_Out),
    .io_MemRLM(_ex2mem_io_MemRLM),
    .io_RtM(_ex2mem_io_RtM),
    .io_BranchJump_JrM(_ex2mem_io_BranchJump_JrM),
    .io_Tlb_ControlM(_ex2mem_io_Tlb_ControlM),
    .io_eBreakM(_ex2mem_io_eBreakM),
    .io_Pc_NextM(_ex2mem_io_Pc_NextM),
    .io_mem_trace_budleM_pc(_ex2mem_io_mem_trace_budleM_pc),
    .io_mem_trace_budleM_data(_ex2mem_io_mem_trace_budleM_data),
    .io_mem_trace_budleM_mem_fetch_type(_ex2mem_io_mem_trace_budleM_mem_fetch_type),
    .io_mem_trace_budleM_addr(_ex2mem_io_mem_trace_budleM_addr),
    .io_mem_trace_budleM_len(_ex2mem_io_mem_trace_budleM_len),
    .io_mem_trace_budleM_cache(_ex2mem_io_mem_trace_budleM_cache),
    .io_CsrWritedataM(_ex2mem_io_CsrWritedataM),
    .io_fence_i_controlM(_ex2mem_io_fence_i_controlM)
  );
  ex2mem _mem2mem2 ( // @[myCPU.scala 128:28]
    .clock(_mem2mem2_clock),
    .reset(_mem2mem2_reset),
    .io1_RegWriteE(_mem2mem2_io1_RegWriteE),
    .io1_MemToRegE(_mem2mem2_io1_MemToRegE),
    .io1_LoadUnsignedE(_mem2mem2_io1_LoadUnsignedE),
    .io1_MemWidthE(_mem2mem2_io1_MemWidthE),
    .io1_csrWriteE(_mem2mem2_io1_csrWriteE),
    .io1_WritecsrAddrE(_mem2mem2_io1_WritecsrAddrE),
    .io1_PCE(_mem2mem2_io1_PCE),
    .io1_MemRLE(_mem2mem2_io1_MemRLE),
    .io1_BranchJump_JrE(_mem2mem2_io1_BranchJump_JrE),
    .io1_Tlb_Control(_mem2mem2_io1_Tlb_Control),
    .io1_eBreakE(_mem2mem2_io1_eBreakE),
    .io1_fence_i_control(_mem2mem2_io1_fence_i_control),
    .io_en(_mem2mem2_io_en),
    .io_clr(_mem2mem2_io_clr),
    .io_WriteDataE(_mem2mem2_io_WriteDataE),
    .io_WriteRegE(_mem2mem2_io_WriteRegE),
    .io_PhyAddrE(_mem2mem2_io_PhyAddrE),
    .io_CsrWritedataE(_mem2mem2_io_CsrWritedataE),
    .io_ExceptionTypeE(_mem2mem2_io_ExceptionTypeE),
    .io_RtE(_mem2mem2_io_RtE),
    .io_Pc_NextE(_mem2mem2_io_Pc_NextE),
    .io_mem_trace_budleE_pc(_mem2mem2_io_mem_trace_budleE_pc),
    .io_mem_trace_budleE_data(_mem2mem2_io_mem_trace_budleE_data),
    .io_mem_trace_budleE_mem_fetch_type(_mem2mem2_io_mem_trace_budleE_mem_fetch_type),
    .io_mem_trace_budleE_addr(_mem2mem2_io_mem_trace_budleE_addr),
    .io_mem_trace_budleE_len(_mem2mem2_io_mem_trace_budleE_len),
    .io_mem_trace_budleE_cache(_mem2mem2_io_mem_trace_budleE_cache),
    .io_RegWriteM(_mem2mem2_io_RegWriteM),
    .io_MemToRegM(_mem2mem2_io_MemToRegM),
    .io_WriteDataM(_mem2mem2_io_WriteDataM),
    .io_WriteRegM(_mem2mem2_io_WriteRegM),
    .io_LoadUnsignedM(_mem2mem2_io_LoadUnsignedM),
    .io_MemWidthM(_mem2mem2_io_MemWidthM),
    .io_PhyAddrM(_mem2mem2_io_PhyAddrM),
    .io_csrWriteM(_mem2mem2_io_csrWriteM),
    .io_WritecsrAddrM(_mem2mem2_io_WritecsrAddrM),
    .io_PCM(_mem2mem2_io_PCM),
    .io_ExceptionTypeM_Out(_mem2mem2_io_ExceptionTypeM_Out),
    .io_MemRLM(_mem2mem2_io_MemRLM),
    .io_RtM(_mem2mem2_io_RtM),
    .io_BranchJump_JrM(_mem2mem2_io_BranchJump_JrM),
    .io_Tlb_ControlM(_mem2mem2_io_Tlb_ControlM),
    .io_eBreakM(_mem2mem2_io_eBreakM),
    .io_Pc_NextM(_mem2mem2_io_Pc_NextM),
    .io_mem_trace_budleM_pc(_mem2mem2_io_mem_trace_budleM_pc),
    .io_mem_trace_budleM_data(_mem2mem2_io_mem_trace_budleM_data),
    .io_mem_trace_budleM_mem_fetch_type(_mem2mem2_io_mem_trace_budleM_mem_fetch_type),
    .io_mem_trace_budleM_addr(_mem2mem2_io_mem_trace_budleM_addr),
    .io_mem_trace_budleM_len(_mem2mem2_io_mem_trace_budleM_len),
    .io_mem_trace_budleM_cache(_mem2mem2_io_mem_trace_budleM_cache),
    .io_CsrWritedataM(_mem2mem2_io_CsrWritedataM),
    .io_fence_i_controlM(_mem2mem2_io_fence_i_controlM)
  );
  id2ex _id2ex ( // @[myCPU.scala 130:26]
    .clock(_id2ex_clock),
    .reset(_id2ex_reset),
    .io1_RegWriteD(_id2ex_io1_RegWriteD),
    .io1_MemToRegD(_id2ex_io1_MemToRegD),
    .io1_MemWriteD(_id2ex_io1_MemWriteD),
    .io1_ALUCtrlD(_id2ex_io1_ALUCtrlD),
    .io1_ALUSrcD_0(_id2ex_io1_ALUSrcD_0),
    .io1_ALUSrcD_1(_id2ex_io1_ALUSrcD_1),
    .io1_RegDstD(_id2ex_io1_RegDstD),
    .io1_LinkD(_id2ex_io1_LinkD),
    .io1_csrWriteD(_id2ex_io1_csrWriteD),
    .io1_csrToRegD(_id2ex_io1_csrToRegD),
    .io1_LoadUnsignedD(_id2ex_io1_LoadUnsignedD),
    .io1_MemWidthD(_id2ex_io1_MemWidthD),
    .io1_ebreakD(_id2ex_io1_ebreakD),
    .io1_data_wD(_id2ex_io1_data_wD),
    .io1_muldiv_control(_id2ex_io1_muldiv_control),
    .io1_muldiv_cal(_id2ex_io1_muldiv_cal),
    .io1_alu_cal(_id2ex_io1_alu_cal),
    .io1_csr_control(_id2ex_io1_csr_control),
    .io1_csr_Imm(_id2ex_io1_csr_Imm),
    .io1_fence_i_control(_id2ex_io1_fence_i_control),
    .io2_RegWriteE(_id2ex_io2_RegWriteE),
    .io2_MemToRegE(_id2ex_io2_MemToRegE),
    .io2_MemWriteE(_id2ex_io2_MemWriteE),
    .io2_ALUCtrlE(_id2ex_io2_ALUCtrlE),
    .io2_ALUSrcE_0(_id2ex_io2_ALUSrcE_0),
    .io2_ALUSrcE_1(_id2ex_io2_ALUSrcE_1),
    .io2_RegDstE(_id2ex_io2_RegDstE),
    .io2_LinkE(_id2ex_io2_LinkE),
    .io2_PCPlus4E(_id2ex_io2_PCPlus4E),
    .io2_LoadUnsignedE(_id2ex_io2_LoadUnsignedE),
    .io2_MemWidthE(_id2ex_io2_MemWidthE),
    .io2_csrWriteE(_id2ex_io2_csrWriteE),
    .io2_WritecsrAddrE(_id2ex_io2_WritecsrAddrE),
    .io2_ReadcsrAddrE(_id2ex_io2_ReadcsrAddrE),
    .io2_PCE(_id2ex_io2_PCE),
    .io2_BranchJump_JrE(_id2ex_io2_BranchJump_JrE),
    .io2_eBreakE(_id2ex_io2_eBreakE),
    .io2_fence_i_control(_id2ex_io2_fence_i_control),
    .io_en(_id2ex_io_en),
    .io_clr(_id2ex_io_clr),
    .io_csrToRegE_Out(_id2ex_io_csrToRegE_Out),
    .io_RD1D(_id2ex_io_RD1D),
    .io_RD2D(_id2ex_io_RD2D),
    .io_R2D(_id2ex_io_R2D),
    .io_R1D(_id2ex_io_R1D),
    .io_ImmD(_id2ex_io_ImmD),
    .io_PCPlus4D(_id2ex_io_PCPlus4D),
    .io_WritecsrAddrD(_id2ex_io_WritecsrAddrD),
    .io_ReadcsrAddrD(_id2ex_io_ReadcsrAddrD),
    .io_PCD(_id2ex_io_PCD),
    .io_ExceptionTypeD(_id2ex_io_ExceptionTypeD),
    .io_Pc_NextD(_id2ex_io_Pc_NextD),
    .io_BranchJump_JrD(_id2ex_io_BranchJump_JrD),
    .io_RD1E(_id2ex_io_RD1E),
    .io_RD2E(_id2ex_io_RD2E),
    .io_R2E(_id2ex_io_R2E),
    .io_R1E(_id2ex_io_R1E),
    .io_ImmE(_id2ex_io_ImmE),
    .io_data_wE(_id2ex_io_data_wE),
    .io_Pc_NextE(_id2ex_io_Pc_NextE),
    .io_muldiv_control(_id2ex_io_muldiv_control),
    .io_alu_calE(_id2ex_io_alu_calE),
    .io_muldiv_calE(_id2ex_io_muldiv_calE),
    .io_ExceptionTypeE_Out(_id2ex_io_ExceptionTypeE_Out),
    .io_csr_controlE(_id2ex_io_csr_controlE),
    .io_csr_ImmE(_id2ex_io_csr_ImmE)
  );
  if2id _if2id ( // @[myCPU.scala 131:26]
    .clock(_if2id_clock),
    .reset(_if2id_reset),
    .io_en(_if2id_io_en),
    .io_clr(_if2id_io_clr),
    .io_InstrF(_if2id_io_InstrF),
    .io_PCPlus4F(_if2id_io_PCPlus4F),
    .io_PCF(_if2id_io_PCF),
    .io_ExceptionTypeF(_if2id_io_ExceptionTypeF),
    .io_InstrD(_if2id_io_InstrD),
    .io_PCPlus4D(_if2id_io_PCPlus4D),
    .io_PCD(_if2id_io_PCD),
    .io_ExceptionTypeD_Out(_if2id_io_ExceptionTypeD_Out)
  );
  mem2wb _mem22wb ( // @[myCPU.scala 133:27]
    .clock(_mem22wb_clock),
    .reset(_mem22wb_reset),
    .io_en(_mem22wb_io_en),
    .io_clr(_mem22wb_io_clr),
    .io_RegWriteM(_mem22wb_io_RegWriteM),
    .io_ResultM(_mem22wb_io_ResultM),
    .io_WriteRegM(_mem22wb_io_WriteRegM),
    .io_csrWriteM(_mem22wb_io_csrWriteM),
    .io_WritecsrAddrM(_mem22wb_io_WritecsrAddrM),
    .io_CsrWritedataM(_mem22wb_io_CsrWritedataM),
    .io_PCM(_mem22wb_io_PCM),
    .io_ExceptionTypeM(_mem22wb_io_ExceptionTypeM),
    .io_BranchJump_JrM(_mem22wb_io_BranchJump_JrM),
    .io_eBreakM(_mem22wb_io_eBreakM),
    .io_Pc_NextM(_mem22wb_io_Pc_NextM),
    .io_Mem_trace_budleM_pc(_mem22wb_io_Mem_trace_budleM_pc),
    .io_Mem_trace_budleM_data(_mem22wb_io_Mem_trace_budleM_data),
    .io_Mem_trace_budleM_mem_fetch_type(_mem22wb_io_Mem_trace_budleM_mem_fetch_type),
    .io_Mem_trace_budleM_addr(_mem22wb_io_Mem_trace_budleM_addr),
    .io_Mem_trace_budleM_len(_mem22wb_io_Mem_trace_budleM_len),
    .io_Mem_trace_budleM_cache(_mem22wb_io_Mem_trace_budleM_cache),
    .io_RegWriteW_Out(_mem22wb_io_RegWriteW_Out),
    .io_ResultW(_mem22wb_io_ResultW),
    .io_WriteRegW(_mem22wb_io_WriteRegW),
    .io_csrWriteW(_mem22wb_io_csrWriteW),
    .io_WritecsrAddrW(_mem22wb_io_WritecsrAddrW),
    .io_PCW(_mem22wb_io_PCW),
    .io_ExceptionTypeW_Out(_mem22wb_io_ExceptionTypeW_Out),
    .io_BranchJump_JrW(_mem22wb_io_BranchJump_JrW),
    .io_eBreakW(_mem22wb_io_eBreakW),
    .io_Pc_NextW(_mem22wb_io_Pc_NextW),
    .io_Mem_trace_budleW_pc(_mem22wb_io_Mem_trace_budleW_pc),
    .io_Mem_trace_budleW_data(_mem22wb_io_Mem_trace_budleW_data),
    .io_Mem_trace_budleW_mem_fetch_type(_mem22wb_io_Mem_trace_budleW_mem_fetch_type),
    .io_Mem_trace_budleW_addr(_mem22wb_io_Mem_trace_budleW_addr),
    .io_Mem_trace_budleW_len(_mem22wb_io_Mem_trace_budleW_len),
    .io_Mem_trace_budleW_cache(_mem22wb_io_Mem_trace_budleW_cache),
    .io_CsrWritedataW(_mem22wb_io_CsrWritedataW)
  );
  addr_cal _addr_cal ( // @[myCPU.scala 134:31]
    .io_d_vaddr(_addr_cal_io_d_vaddr),
    .io_d_paddr(_addr_cal_io_d_paddr),
    .io_d_cached(_addr_cal_io_d_cached)
  );
  muldiv _muldiv ( // @[myCPU.scala 135:26]
    .clock(_muldiv_clock),
    .reset(_muldiv_reset),
    .io_en(_muldiv_io_en),
    .io_ctrl(_muldiv_io_ctrl),
    .io_in1(_muldiv_io_in1),
    .io_in2(_muldiv_io_in2),
    .io_data_out(_muldiv_io_data_out),
    .io_pending(_muldiv_io_pending)
  );
  regfile _regfile ( // @[myCPU.scala 137:26]
    .clock(_regfile_clock),
    .reset(_regfile_reset),
    .io_A1(_regfile_io_A1),
    .io_A2(_regfile_io_A2),
    .io_WE3(_regfile_io_WE3),
    .io_A3(_regfile_io_A3),
    .io_WD3(_regfile_io_WD3),
    .io_RD1(_regfile_io_RD1),
    .io_RD2(_regfile_io_RD2),
    .io_reg_file_alL_out(_regfile_io_reg_file_alL_out)
  );
  mem_trace_module _mtrace_mod ( // @[myCPU.scala 138:29]
    .reset(_mtrace_mod_reset),
    .clock(_mtrace_mod_clock),
    .data(_mtrace_mod_data),
    .pc(_mtrace_mod_pc),
    .addr(_mtrace_mod_addr),
    .mem_req(_mtrace_mod_mem_req),
    .mem_write_read(_mtrace_mod_mem_write_read),
    .mem_size(_mtrace_mod_mem_size),
    .mem_cached(_mtrace_mod_mem_cached)
  );
  fifo_with_bundle fifo_with_bundle ( // @[myCPU.scala 159:29]
    .clock(fifo_with_bundle_clock),
    .reset(fifo_with_bundle_reset),
    .io_read_en(fifo_with_bundle_io_read_en),
    .io_write_en(fifo_with_bundle_io_write_en),
    .io_read_out_0_pc(fifo_with_bundle_io_read_out_0_pc),
    .io_read_out_0_inst(fifo_with_bundle_io_read_out_0_inst),
    .io_read_out_0_exception_type(fifo_with_bundle_io_read_out_0_exception_type),
    .io_read_out_0_pre_pc_target(fifo_with_bundle_io_read_out_0_pre_pc_target),
    .io_read_out_0_pre_lookup_data(fifo_with_bundle_io_read_out_0_pre_lookup_data),
    .io_read_out_0_pre_hashcode(fifo_with_bundle_io_read_out_0_pre_hashcode),
    .io_read_out_0_pre_pht(fifo_with_bundle_io_read_out_0_pre_pht),
    .io_read_out_0_pre_bht(fifo_with_bundle_io_read_out_0_pre_bht),
    .io_read_out_0_pre_lookup_value(fifo_with_bundle_io_read_out_0_pre_lookup_value),
    .io_read_out_0_pre_decoder_branchD_flag(fifo_with_bundle_io_read_out_0_pre_decoder_branchD_flag),
    .io_read_out_0_pre_decoder_jump(fifo_with_bundle_io_read_out_0_pre_decoder_jump),
    .io_read_out_0_pre_decoder_branchdata(fifo_with_bundle_io_read_out_0_pre_decoder_branchdata),
    .io_read_out_0_pre_decoder_jr(fifo_with_bundle_io_read_out_0_pre_decoder_jr),
    .io_read_out_0_true_branch_state(fifo_with_bundle_io_read_out_0_true_branch_state),
    .io_write_in_0_pc(fifo_with_bundle_io_write_in_0_pc),
    .io_write_in_0_inst(fifo_with_bundle_io_write_in_0_inst),
    .io_write_in_0_pre_pc_target(fifo_with_bundle_io_write_in_0_pre_pc_target),
    .io_write_in_0_pre_lookup_data(fifo_with_bundle_io_write_in_0_pre_lookup_data),
    .io_write_in_0_pre_hashcode(fifo_with_bundle_io_write_in_0_pre_hashcode),
    .io_write_in_0_pre_pht(fifo_with_bundle_io_write_in_0_pre_pht),
    .io_write_in_0_pre_bht(fifo_with_bundle_io_write_in_0_pre_bht),
    .io_write_in_0_pre_lookup_value(fifo_with_bundle_io_write_in_0_pre_lookup_value),
    .io_write_in_0_pre_decoder_branchD_flag(fifo_with_bundle_io_write_in_0_pre_decoder_branchD_flag),
    .io_write_in_0_pre_decoder_jump(fifo_with_bundle_io_write_in_0_pre_decoder_jump),
    .io_write_in_0_pre_decoder_branchdata(fifo_with_bundle_io_write_in_0_pre_decoder_branchdata),
    .io_write_in_0_pre_decoder_jr(fifo_with_bundle_io_write_in_0_pre_decoder_jr),
    .io_write_in_0_true_branch_state(fifo_with_bundle_io_write_in_0_true_branch_state),
    .io_full(fifo_with_bundle_io_full),
    .io_empty(fifo_with_bundle_io_empty),
    .io_point_write_en(fifo_with_bundle_io_point_write_en),
    .io_point_flush(fifo_with_bundle_io_point_flush)
  );
  pc_detail stage_fec_1_pc_L ( // @[myCPU.scala 421:34]
    .clock(stage_fec_1_pc_L_clock),
    .reset(stage_fec_1_pc_L_reset),
    .io_stall(stage_fec_1_pc_L_io_stall),
    .io_flush(stage_fec_1_pc_L_io_flush),
    .io_in_pc_value_in(stage_fec_1_pc_L_io_in_pc_value_in),
    .io_out_pc_value_out(stage_fec_1_pc_L_io_out_pc_value_out)
  );
  pc_detail stage_fec_1_pc_M ( // @[myCPU.scala 422:34]
    .clock(stage_fec_1_pc_M_clock),
    .reset(stage_fec_1_pc_M_reset),
    .io_stall(stage_fec_1_pc_M_io_stall),
    .io_flush(stage_fec_1_pc_M_io_flush),
    .io_in_pc_value_in(stage_fec_1_pc_M_io_in_pc_value_in),
    .io_out_pc_value_out(stage_fec_1_pc_M_io_out_pc_value_out)
  );
  pc_detail stage_fec_1_pc_R ( // @[myCPU.scala 423:34]
    .clock(stage_fec_1_pc_R_clock),
    .reset(stage_fec_1_pc_R_reset),
    .io_stall(stage_fec_1_pc_R_io_stall),
    .io_flush(stage_fec_1_pc_R_io_flush),
    .io_in_pc_value_in(stage_fec_1_pc_R_io_in_pc_value_in),
    .io_out_pc_value_out(stage_fec_1_pc_R_io_out_pc_value_out)
  );
  branch_prediction_with_blockram branch_prediction_with_blockram ( // @[myCPU.scala 452:21]
    .clock(branch_prediction_with_blockram_clock),
    .reset(branch_prediction_with_blockram_reset),
    .io_pc(branch_prediction_with_blockram_io_pc),
    .io_write_pc(branch_prediction_with_blockram_io_write_pc),
    .io_aw_pht_ways_addr(branch_prediction_with_blockram_io_aw_pht_ways_addr),
    .io_aw_pht_addr(branch_prediction_with_blockram_io_aw_pht_addr),
    .io_aw_bht_addr(branch_prediction_with_blockram_io_aw_bht_addr),
    .io_aw_target_addr(branch_prediction_with_blockram_io_aw_target_addr),
    .io_btb_write(branch_prediction_with_blockram_io_btb_write),
    .io_bht_write(branch_prediction_with_blockram_io_bht_write),
    .io_pht_write(branch_prediction_with_blockram_io_pht_write),
    .io_bht_in(branch_prediction_with_blockram_io_bht_in),
    .io_pht_in(branch_prediction_with_blockram_io_pht_in),
    .io_out_L(branch_prediction_with_blockram_io_out_L),
    .io_pre_L(branch_prediction_with_blockram_io_pre_L),
    .io_bht_L(branch_prediction_with_blockram_io_bht_L),
    .io_btb_hit_0(branch_prediction_with_blockram_io_btb_hit_0),
    .io_pre_target_L(branch_prediction_with_blockram_io_pre_target_L),
    .io_stage2_stall(branch_prediction_with_blockram_io_stage2_stall),
    .io_stage2_flush(branch_prediction_with_blockram_io_stage2_flush),
    .io_pht_lookup_value_out(branch_prediction_with_blockram_io_pht_lookup_value_out),
    .io_lookup_data_0(branch_prediction_with_blockram_io_lookup_data_0)
  );
  pc_detail stage_fec_2_pc_L ( // @[myCPU.scala 521:34]
    .clock(stage_fec_2_pc_L_clock),
    .reset(stage_fec_2_pc_L_reset),
    .io_stall(stage_fec_2_pc_L_io_stall),
    .io_flush(stage_fec_2_pc_L_io_flush),
    .io_in_pc_value_in(stage_fec_2_pc_L_io_in_pc_value_in),
    .io_out_pc_value_out(stage_fec_2_pc_L_io_out_pc_value_out)
  );
  pc_detail stage_fec_2_pc_M ( // @[myCPU.scala 522:34]
    .clock(stage_fec_2_pc_M_clock),
    .reset(stage_fec_2_pc_M_reset),
    .io_stall(stage_fec_2_pc_M_io_stall),
    .io_flush(stage_fec_2_pc_M_io_flush),
    .io_in_pc_value_in(stage_fec_2_pc_M_io_in_pc_value_in),
    .io_out_pc_value_out(stage_fec_2_pc_M_io_out_pc_value_out)
  );
  pc_detail stage_fec_2_pc_R ( // @[myCPU.scala 523:34]
    .clock(stage_fec_2_pc_R_clock),
    .reset(stage_fec_2_pc_R_reset),
    .io_stall(stage_fec_2_pc_R_io_stall),
    .io_flush(stage_fec_2_pc_R_io_flush),
    .io_in_pc_value_in(stage_fec_2_pc_R_io_in_pc_value_in),
    .io_out_pc_value_out(stage_fec_2_pc_R_io_out_pc_value_out)
  );
  bru_detail id_bru_state ( // @[myCPU.scala 685:31]
    .clock(id_bru_state_clock),
    .reset(id_bru_state_reset),
    .io_stall(id_bru_state_io_stall),
    .io_flush(id_bru_state_io_flush),
    .io_in_pht(id_bru_state_io_in_pht),
    .io_in_bht(id_bru_state_io_in_bht),
    .io_in_hashcode(id_bru_state_io_in_hashcode),
    .io_in_target_pc(id_bru_state_io_in_target_pc),
    .io_in_lookup_data(id_bru_state_io_in_lookup_data),
    .io_in_pht_lookup_value(id_bru_state_io_in_pht_lookup_value),
    .io_out_pht(id_bru_state_io_out_pht),
    .io_out_bht(id_bru_state_io_out_bht),
    .io_out_hashcode(id_bru_state_io_out_hashcode),
    .io_out_target_pc(id_bru_state_io_out_target_pc),
    .io_out_lookup_data(id_bru_state_io_out_lookup_data),
    .io_out_pht_lookup_value(id_bru_state_io_out_pht_lookup_value)
  );
  bru_detail ex_bru_state ( // @[myCPU.scala 689:31]
    .clock(ex_bru_state_clock),
    .reset(ex_bru_state_reset),
    .io_stall(ex_bru_state_io_stall),
    .io_flush(ex_bru_state_io_flush),
    .io_in_pht(ex_bru_state_io_in_pht),
    .io_in_bht(ex_bru_state_io_in_bht),
    .io_in_hashcode(ex_bru_state_io_in_hashcode),
    .io_in_target_pc(ex_bru_state_io_in_target_pc),
    .io_in_lookup_data(ex_bru_state_io_in_lookup_data),
    .io_in_pht_lookup_value(ex_bru_state_io_in_pht_lookup_value),
    .io_out_pht(ex_bru_state_io_out_pht),
    .io_out_bht(ex_bru_state_io_out_bht),
    .io_out_hashcode(ex_bru_state_io_out_hashcode),
    .io_out_target_pc(ex_bru_state_io_out_target_pc),
    .io_out_lookup_data(ex_bru_state_io_out_lookup_data),
    .io_out_pht_lookup_value(ex_bru_state_io_out_pht_lookup_value)
  );
  bru_detail mem_bru_state ( // @[myCPU.scala 693:32]
    .clock(mem_bru_state_clock),
    .reset(mem_bru_state_reset),
    .io_stall(mem_bru_state_io_stall),
    .io_flush(mem_bru_state_io_flush),
    .io_in_pht(mem_bru_state_io_in_pht),
    .io_in_bht(mem_bru_state_io_in_bht),
    .io_in_hashcode(mem_bru_state_io_in_hashcode),
    .io_in_target_pc(mem_bru_state_io_in_target_pc),
    .io_in_lookup_data(mem_bru_state_io_in_lookup_data),
    .io_in_pht_lookup_value(mem_bru_state_io_in_pht_lookup_value),
    .io_out_pht(mem_bru_state_io_out_pht),
    .io_out_bht(mem_bru_state_io_out_bht),
    .io_out_hashcode(mem_bru_state_io_out_hashcode),
    .io_out_target_pc(mem_bru_state_io_out_target_pc),
    .io_out_lookup_data(mem_bru_state_io_out_lookup_data),
    .io_out_pht_lookup_value(mem_bru_state_io_out_pht_lookup_value)
  );
  bru_detail mem2_bru_state ( // @[myCPU.scala 697:33]
    .clock(mem2_bru_state_clock),
    .reset(mem2_bru_state_reset),
    .io_stall(mem2_bru_state_io_stall),
    .io_flush(mem2_bru_state_io_flush),
    .io_in_pht(mem2_bru_state_io_in_pht),
    .io_in_bht(mem2_bru_state_io_in_bht),
    .io_in_hashcode(mem2_bru_state_io_in_hashcode),
    .io_in_target_pc(mem2_bru_state_io_in_target_pc),
    .io_in_lookup_data(mem2_bru_state_io_in_lookup_data),
    .io_in_pht_lookup_value(mem2_bru_state_io_in_pht_lookup_value),
    .io_out_pht(mem2_bru_state_io_out_pht),
    .io_out_bht(mem2_bru_state_io_out_bht),
    .io_out_hashcode(mem2_bru_state_io_out_hashcode),
    .io_out_target_pc(mem2_bru_state_io_out_target_pc),
    .io_out_lookup_data(mem2_bru_state_io_out_lookup_data),
    .io_out_pht_lookup_value(mem2_bru_state_io_out_pht_lookup_value)
  );
  bru_detail wb_bru_state ( // @[myCPU.scala 701:31]
    .clock(wb_bru_state_clock),
    .reset(wb_bru_state_reset),
    .io_stall(wb_bru_state_io_stall),
    .io_flush(wb_bru_state_io_flush),
    .io_in_pht(wb_bru_state_io_in_pht),
    .io_in_bht(wb_bru_state_io_in_bht),
    .io_in_hashcode(wb_bru_state_io_in_hashcode),
    .io_in_target_pc(wb_bru_state_io_in_target_pc),
    .io_in_lookup_data(wb_bru_state_io_in_lookup_data),
    .io_in_pht_lookup_value(wb_bru_state_io_in_pht_lookup_value),
    .io_out_pht(wb_bru_state_io_out_pht),
    .io_out_bht(wb_bru_state_io_out_bht),
    .io_out_hashcode(wb_bru_state_io_out_hashcode),
    .io_out_target_pc(wb_bru_state_io_out_target_pc),
    .io_out_lookup_data(wb_bru_state_io_out_lookup_data),
    .io_out_pht_lookup_value(wb_bru_state_io_out_pht_lookup_value)
  );
  difftest_commit _commit_difftest ( // @[myCPU.scala 1148:34]
    .reset(_commit_difftest_reset),
    .clock(_commit_difftest_clock),
    .gpr_wire(_commit_difftest_gpr_wire),
    .pc(_commit_difftest_pc),
    .debug_pc(_commit_difftest_debug_pc),
    .inst_commit(_commit_difftest_inst_commit),
    .data_ok_ok(_commit_difftest_data_ok_ok),
    .cpu_ebreak_sign(_commit_difftest_cpu_ebreak_sign)
  );
  assign inst_cache = Pc_Next[31:29] == 3'h4; // @[macros.scala 479:55]
  assign inst_sram_en = stage2_stall; // @[myCPU.scala 384:17]
  assign inst_sram_addr = _stage_fec_2_branch_answer_T_7 ? _csr_io_return_pc : _Pc_Next_T_3; // @[myCPU.scala 377:19]
  assign stage2_flush = fifo_with_bundle_io_point_write_en & _stage_fec_2_data_valid_T | _stage_fec_2_branch_answer_T_7; // @[myCPU.scala 581:72]
  assign stage1_valid_flush = _pc_next_wait_T | _stage_fec_2_branch_answer_T_7; // @[myCPU.scala 591:85]
  assign inst_ready_to_use = Pc_Next[1:0] == 2'h0; // @[myCPU.scala 385:39]
  assign inst_buffer_full = fifo_with_bundle_io_full; // @[myCPU.scala 600:22]
  assign data_sram_en = _dmemreq_io_req & ~_dmem_io_data_pending; // @[myCPU.scala 239:44]
  assign data_sram_wen = _dmemreq_io_wr; // @[myCPU.scala 245:13]
  assign data_size = _dmemreq_io_size; // @[myCPU.scala 1205:15]
  assign data_sram_addr = _dmemreq_io_addr; // @[myCPU.scala 241:15]
  assign data_sram_wdata = _dmemreq_io_wdata; // @[myCPU.scala 242:16]
  assign data_cache = _addr_cal_io_d_cached; // @[myCPU.scala 1204:63]
  assign data_wstrb = _dmemreq_io_wstrb; // @[myCPU.scala 243:16]
  assign data_fence_i_control = _ex2mem_io_fence_i_controlM; // @[myCPU.scala 954:26]
  assign debug_wb_pc = _mem22wb_io_PCW; // @[myCPU.scala 303:17]
  assign debug_wb_rf_wen = reg_pc == _mem22wb_io_PCW ? 4'h0 : _debug_wb_rf_wen_T_2; // @[myCPU.scala 304:27]
  assign debug_wb_rf_wnum = _regfile_io_A3; // @[myCPU.scala 305:22]
  assign debug_wb_rf_wdata = _regfile_io_WD3; // @[myCPU.scala 306:23]
  assign icache_tag_flush = _csr_io_icache_tags_flush; // @[myCPU.scala 1215:22]
  assign _alu_io_ctrl = _id2ex_io2_ALUCtrlE; // @[myCPU.scala 891:18]
  assign _alu_io_in1 = {Src1E[63:32],Src1E[31:0]}; // @[Cat.scala 31:58]
  assign _alu_io_in2 = {Src2E[63:32],Src2E[31:0]}; // @[Cat.scala 31:58]
  assign _alu_io_data_w = _id2ex_io_data_wE; // @[myCPU.scala 892:20]
  assign _br_reset = ~resetn; // @[myCPU.scala 114:41]
  assign _br_io_r1 = _cfu_io_Forward1D[0] ? resultE2M_Reg : _BranchR1D_T_2; // @[myCPU.scala 773:20]
  assign _br_io_r2 = _cfu_io_Forward2D[0] ? resultE2M_Reg : _BranchR2D_T_2; // @[myCPU.scala 775:20]
  assign _br_io_branch = pre_decoder_branchdata; // @[myCPU.scala 783:19]
  assign _cfu_reset = ~resetn; // @[myCPU.scala 114:41]
  assign _cfu_io_Inst_Fifo_Empty = fifo_with_bundle_io_empty; // @[myCPU.scala 584:29]
  assign _cfu_io_dmem_calD = _cu_io1_dmem_addr_cal; // @[myCPU.scala 835:23]
  assign _cfu_io_BranchD_Flag = pre_decoder_branchD_flag; // @[myCPU.scala 1237:26]
  assign _cfu_io_JRD = pre_decoder_jr; // @[myCPU.scala 1233:25]
  assign _cfu_io_CanBranchD = ~(id_exception | ex_exception | mem_exception | mem2_exception | wb_exception); // @[myCPU.scala 1234:111]
  assign _cfu_io_DivPendingE = _muldiv_io_pending; // @[myCPU.scala 1238:33]
  assign _cfu_io_DataPendingM = _dmem_io_data_pending; // @[myCPU.scala 1240:33]
  assign _cfu_io_InException = _csr_io_exception; // @[myCPU.scala 1227:25]
  assign _cfu_io_WriteRegE = _id2ex_io2_RegDstE; // @[myCPU.scala 1244:33]
  assign _cfu_io_RegWriteE = _id2ex_io2_RegWriteE; // @[myCPU.scala 1246:33]
  assign _cfu_io_csrToRegE = _id2ex_io_ExceptionTypeE_Out == 32'h0 & _id2ex_io_csrToRegE_Out; // @[myCPU.scala 887:24]
  assign _cfu_io_WriteRegM = _ex2mem_io_WriteRegM; // @[myCPU.scala 1250:33]
  assign _cfu_io_MemToRegM = _ex2mem_io_MemToRegM; // @[myCPU.scala 1251:33]
  assign _cfu_io_RegWriteM = _ex2mem_io_RegWriteM; // @[myCPU.scala 1252:33]
  assign _cfu_io_csrWriteM = _ex2mem_io_csrWriteM; // @[myCPU.scala 1253:33]
  assign _cfu_io_WriteRegM2 = _mem2mem2_io_WriteRegM; // @[myCPU.scala 1274:25]
  assign _cfu_io_MemToRegM2 = _mem2mem2_io_MemToRegM; // @[myCPU.scala 1275:25]
  assign _cfu_io_RegWriteM2 = _mem2mem2_io_RegWriteM; // @[myCPU.scala 1276:25]
  assign _cfu_io_csrWriteM2 = _mem2mem2_io_csrWriteM; // @[myCPU.scala 1272:24]
  assign _cfu_io_WriteRegW = _mem22wb_io_WriteRegW; // @[myCPU.scala 1263:33]
  assign _cfu_io_RegWriteW = wb_exception ? 1'h0 : _mem22wb_io_RegWriteW_Out; // @[myCPU.scala 1162:21]
  assign _cfu_io_ReadcsrAddrE = _id2ex_io2_ReadcsrAddrE; // @[myCPU.scala 1255:34]
  assign _cfu_io_WritecsrAddrM = _ex2mem_io_WritecsrAddrM; // @[myCPU.scala 1258:34]
  assign _cfu_io_WritecsrAddrM2 = _mem2mem2_io_WritecsrAddrM; // @[myCPU.scala 1273:28]
  assign _cfu_io_R2D = _if2id_io_InstrD[24:20]; // @[myCPU.scala 205:27]
  assign _cfu_io_R1D = _if2id_io_InstrD[19:15]; // @[myCPU.scala 206:27]
  assign _cfu_io_R2E = _id2ex_io_R2E; // @[myCPU.scala 1269:33]
  assign _cfu_io_R1E = _id2ex_io_R1E; // @[myCPU.scala 1268:33]
  assign _csr_clock = clk; // @[myCPU.scala 114:23]
  assign _csr_reset = ~resetn; // @[myCPU.scala 114:41]
  assign _csr_io_csr_read_addr = _id2ex_io2_ReadcsrAddrE; // @[myCPU.scala 970:27]
  assign _csr_io_csr_write_addr = _mem22wb_io_WritecsrAddrW; // @[myCPU.scala 971:28]
  assign _csr_io_csr_write_data = _mem22wb_io_CsrWritedataW; // @[myCPU.scala 1222:30]
  assign _csr_io_csr_write_en = csrWriteW | tlb_exception_co0_writeW; // @[myCPU.scala 1212:47]
  assign _csr_io_pc = _PCW_Reg_T ? _mem22wb_io_PCW : PCW_Reg; // @[myCPU.scala 1210:25]
  assign _csr_io_exception_type_i = _mem22wb_io_ExceptionTypeW_Out; // @[myCPU.scala 1213:30]
  assign _csr_io_int_type_timer = int_instanceW_timer; // @[myCPU.scala 1209:22]
  assign _cu_io1_InstrD = _if2id_io_InstrD; // @[myCPU.scala 771:20]
  assign _dmem_io_data_ok = data_stage2_stall; // @[myCPU.scala 266:25]
  assign _dmem_io_rdata = data_sram_rdata; // @[myCPU.scala 267:25]
  assign _dmem_io_Physisc_Address = _mem2mem2_io_PhyAddrM; // @[myCPU.scala 271:30]
  assign _dmem_io_WIDTH = _mem2mem2_io_MemWidthM; // @[myCPU.scala 269:25]
  assign _dmem_io_SIGN = ~_mem2mem2_io_LoadUnsignedM; // @[myCPU.scala 270:22]
  assign _dmemreq_io_en = _T_37 ? 1'h0 : _commit_cache_reg_T; // @[myCPU.scala 909:26]
  assign _dmemreq_io_MemWriteE = _id2ex_io2_MemWriteE; // @[myCPU.scala 915:27]
  assign _dmemreq_io_MemToRegE = _id2ex_io2_MemToRegE; // @[myCPU.scala 912:27]
  assign _dmemreq_io_MemWidthE = _id2ex_io2_MemWidthE; // @[myCPU.scala 913:27]
  assign _dmemreq_io_VAddrE = _addr_cal_io_d_paddr; // @[myCPU.scala 1199:23]
  assign _dmemreq_io_WriteDataE = Forward_Lock2E ? RD2ForWardE_r : RD2ForWardE_p; // @[myCPU.scala 855:23]
  assign _ex2mem_clock = clk; // @[myCPU.scala 114:23]
  assign _ex2mem_reset = ~resetn; // @[myCPU.scala 114:41]
  assign _ex2mem_io1_RegWriteE = _id2ex_io2_RegWriteE; // @[myCPU.scala 165:15]
  assign _ex2mem_io1_MemToRegE = _id2ex_io2_MemToRegE; // @[myCPU.scala 165:15]
  assign _ex2mem_io1_LoadUnsignedE = _id2ex_io2_LoadUnsignedE; // @[myCPU.scala 165:15]
  assign _ex2mem_io1_MemWidthE = _id2ex_io2_MemWidthE; // @[myCPU.scala 165:15]
  assign _ex2mem_io1_csrWriteE = _id2ex_io2_csrWriteE; // @[myCPU.scala 165:15]
  assign _ex2mem_io1_WritecsrAddrE = _id2ex_io2_WritecsrAddrE; // @[myCPU.scala 165:15]
  assign _ex2mem_io1_PCE = _id2ex_io2_PCE; // @[myCPU.scala 165:15]
  assign _ex2mem_io1_MemRLE = 2'h0; // @[myCPU.scala 165:15]
  assign _ex2mem_io1_BranchJump_JrE = _id2ex_io2_BranchJump_JrE; // @[myCPU.scala 165:15]
  assign _ex2mem_io1_Tlb_Control = 3'h0; // @[myCPU.scala 165:15]
  assign _ex2mem_io1_eBreakE = _id2ex_io2_eBreakE; // @[myCPU.scala 165:15]
  assign _ex2mem_io1_fence_i_control = _id2ex_io2_fence_i_control; // @[myCPU.scala 165:15]
  assign _ex2mem_io_en = _cfu_io_StallE; // @[myCPU.scala 212:30]
  assign _ex2mem_io_clr = _cfu_io_FlushM; // @[myCPU.scala 213:30]
  assign _ex2mem_io_WriteDataE = Forward_Lock2E ? RD2ForWardE_r : RD2ForWardE_p; // @[myCPU.scala 855:23]
  assign _ex2mem_io_WriteRegE = _id2ex_io2_RegDstE; // @[myCPU.scala 942:26]
  assign _ex2mem_io_PhyAddrE = _addr_cal_io_d_paddr; // @[myCPU.scala 945:27]
  assign _ex2mem_io_CsrWritedataE = _CalCsrDataE_T_12 | _CalCsrDataE_T_11; // @[Mux.scala 27:73]
  assign _ex2mem_io_ExceptionTypeE = _id2ex_io_ExceptionTypeE_Out != 32'h0 ? _id2ex_io_ExceptionTypeE_Out : {{19'd0},
    _temp_exceptionE_T_11}; // @[myCPU.scala 926:30]
  assign _ex2mem_io_RtE = Forward_Lock2E ? RD2ForWardE_r : RD2ForWardE_p; // @[myCPU.scala 855:23]
  assign _ex2mem_io_Pc_NextE = _id2ex_io_Pc_NextE; // @[myCPU.scala 934:25]
  assign _ex2mem_io_mem_trace_budleE_pc = _id2ex_io2_PCE; // @[myCPU.scala 947:36]
  assign _ex2mem_io_mem_trace_budleE_data = data_sram_wdata; // @[myCPU.scala 948:38]
  assign _ex2mem_io_mem_trace_budleE_mem_fetch_type = {_id2ex_io2_MemToRegE,_id2ex_io2_MemWriteE}; // @[Cat.scala 31:58]
  assign _ex2mem_io_mem_trace_budleE_addr = data_sram_addr; // @[myCPU.scala 950:48]
  assign _ex2mem_io_mem_trace_budleE_len = {{1'd0}, data_size}; // @[myCPU.scala 951:48]
  assign _ex2mem_io_mem_trace_budleE_cache = data_cache; // @[myCPU.scala 952:48]
  assign _mem2mem2_clock = clk; // @[myCPU.scala 114:23]
  assign _mem2mem2_reset = ~resetn; // @[myCPU.scala 114:41]
  assign _mem2mem2_io1_RegWriteE = _ex2mem_io_RegWriteM; // @[myCPU.scala 1057:30]
  assign _mem2mem2_io1_MemToRegE = _ex2mem_io_MemToRegM; // @[myCPU.scala 1058:30]
  assign _mem2mem2_io1_LoadUnsignedE = _ex2mem_io_LoadUnsignedM; // @[myCPU.scala 1062:30]
  assign _mem2mem2_io1_MemWidthE = _ex2mem_io_MemWidthM; // @[myCPU.scala 1063:30]
  assign _mem2mem2_io1_csrWriteE = __mem2mem2_io_csrWriteE_T | _ex2mem_io_Tlb_ControlM[2]; // @[myCPU.scala 1066:61]
  assign _mem2mem2_io1_WritecsrAddrE = inst_tlb_exceptionM ? 12'ha : _ex2mem_io_WritecsrAddrM; // @[myCPU.scala 1067:36]
  assign _mem2mem2_io1_PCE = _ex2mem_io_PCM; // @[myCPU.scala 1068:30]
  assign _mem2mem2_io1_MemRLE = _ex2mem_io_MemRLM; // @[myCPU.scala 1070:30]
  assign _mem2mem2_io1_BranchJump_JrE = _ex2mem_io_BranchJump_JrM; // @[myCPU.scala 1071:30]
  assign _mem2mem2_io1_Tlb_Control = _ex2mem_io_Tlb_ControlM; // @[myCPU.scala 1080:27]
  assign _mem2mem2_io1_eBreakE = _ex2mem_io1_eBreakE; // @[myCPU.scala 1045:24]
  assign _mem2mem2_io1_fence_i_control = _ex2mem_io_fence_i_controlM; // @[myCPU.scala 1055:31]
  assign _mem2mem2_io_en = _cfu_io_StallM2; // @[myCPU.scala 1099:20]
  assign _mem2mem2_io_clr = _cfu_io_FlushM2; // @[myCPU.scala 1098:20]
  assign _mem2mem2_io_WriteDataE = _ex2mem_io_WriteDataM; // @[myCPU.scala 1095:30]
  assign _mem2mem2_io_WriteRegE = _ex2mem_io_WriteRegM; // @[myCPU.scala 1046:24]
  assign _mem2mem2_io_PhyAddrE = _ex2mem_io_PhyAddrM; // @[myCPU.scala 1047:23]
  assign _mem2mem2_io_CsrWritedataE = _ex2mem_io_CsrWritedataM; // @[myCPU.scala 1081:29]
  assign _mem2mem2_io_ExceptionTypeE = mem_exception ? _ex2mem_io_ExceptionTypeM_Out : 32'h0; // @[myCPU.scala 1039:21]
  assign _mem2mem2_io_RtE = _ex2mem_io_RtM; // @[myCPU.scala 1053:18]
  assign _mem2mem2_io_Pc_NextE = _ex2mem_io_Pc_NextM; // @[myCPU.scala 1044:24]
  assign _mem2mem2_io_mem_trace_budleE_pc = _ex2mem_io_mem_trace_budleM_pc; // @[myCPU.scala 1054:31]
  assign _mem2mem2_io_mem_trace_budleE_data = _ex2mem_io_mem_trace_budleM_data; // @[myCPU.scala 1054:31]
  assign _mem2mem2_io_mem_trace_budleE_mem_fetch_type = _ex2mem_io_mem_trace_budleM_mem_fetch_type; // @[myCPU.scala 1054:31]
  assign _mem2mem2_io_mem_trace_budleE_addr = _ex2mem_io_mem_trace_budleM_addr; // @[myCPU.scala 1054:31]
  assign _mem2mem2_io_mem_trace_budleE_len = _ex2mem_io_mem_trace_budleM_len; // @[myCPU.scala 1054:31]
  assign _mem2mem2_io_mem_trace_budleE_cache = _ex2mem_io_mem_trace_budleM_cache; // @[myCPU.scala 1054:31]
  assign _id2ex_clock = clk; // @[myCPU.scala 114:23]
  assign _id2ex_reset = ~resetn; // @[myCPU.scala 114:41]
  assign _id2ex_io1_RegWriteD = _cu_io_RegWriteD; // @[myCPU.scala 164:15]
  assign _id2ex_io1_MemToRegD = _cu_io_MemToRegD; // @[myCPU.scala 164:15]
  assign _id2ex_io1_MemWriteD = _cu_io_MemWriteD; // @[myCPU.scala 164:15]
  assign _id2ex_io1_ALUCtrlD = _cu_io_ALUCtrlD; // @[myCPU.scala 164:15]
  assign _id2ex_io1_ALUSrcD_0 = _cu_io_ALUSrcD_0; // @[myCPU.scala 164:15]
  assign _id2ex_io1_ALUSrcD_1 = _cu_io_ALUSrcD_1; // @[myCPU.scala 164:15]
  assign _id2ex_io1_RegDstD = _cu_io_RegDstD; // @[myCPU.scala 164:15]
  assign _id2ex_io1_LinkD = _cu_io_LinkD; // @[myCPU.scala 164:15]
  assign _id2ex_io1_csrWriteD = _cu_io_csrWriteD; // @[myCPU.scala 164:15]
  assign _id2ex_io1_csrToRegD = _cu_io_csrToRegD; // @[myCPU.scala 164:15]
  assign _id2ex_io1_LoadUnsignedD = _cu_io_LoadUnsignedD; // @[myCPU.scala 164:15]
  assign _id2ex_io1_MemWidthD = _cu_io_MemWidthD; // @[myCPU.scala 164:15]
  assign _id2ex_io1_ebreakD = _cu_io_ebreakD; // @[myCPU.scala 164:15]
  assign _id2ex_io1_data_wD = _cu_io_data_wD; // @[myCPU.scala 164:15]
  assign _id2ex_io1_muldiv_control = _cu_io_muldiv_control; // @[myCPU.scala 164:15]
  assign _id2ex_io1_muldiv_cal = _cu_io_muldiv_cal; // @[myCPU.scala 164:15]
  assign _id2ex_io1_alu_cal = _cu_io_alu_cal; // @[myCPU.scala 164:15]
  assign _id2ex_io1_csr_control = _cu_io_csr_control; // @[myCPU.scala 164:15]
  assign _id2ex_io1_csr_Imm = _cu_io_csr_Imm; // @[myCPU.scala 164:15]
  assign _id2ex_io1_fence_i_control = _cu_io_fence_i_control; // @[myCPU.scala 164:15]
  assign _id2ex_io_en = _cfu_io_StallD; // @[myCPU.scala 193:29]
  assign _id2ex_io_clr = _cfu_io_FlushE; // @[myCPU.scala 194:29]
  assign _id2ex_io_RD1D = _cfu_io_Forward1D[0] ? resultE2M_Reg : _BranchR1D_T_2; // @[myCPU.scala 813:25]
  assign _id2ex_io_RD2D = _cfu_io_Forward2D[0] ? resultE2M_Reg : _BranchR2D_T_2; // @[myCPU.scala 814:25]
  assign _id2ex_io_R2D = _if2id_io_InstrD[24:20]; // @[myCPU.scala 205:27]
  assign _id2ex_io_R1D = _if2id_io_InstrD[19:15]; // @[myCPU.scala 206:27]
  assign _id2ex_io_ImmD = _cu_io_ImmD; // @[myCPU.scala 812:19]
  assign _id2ex_io_PCPlus4D = _if2id_io_PCPlus4D; // @[myCPU.scala 825:29]
  assign _id2ex_io_WritecsrAddrD = _if2id_io_InstrD[31:20]; // @[myCPU.scala 815:38]
  assign _id2ex_io_ReadcsrAddrD = _if2id_io_InstrD[31:20]; // @[myCPU.scala 817:38]
  assign _id2ex_io_PCD = _if2id_io_PCD; // @[myCPU.scala 826:28]
  assign _id2ex_io_ExceptionTypeD = __id2ex_io_ExceptionTypeD_T_13[31:0]; // @[myCPU.scala 802:31]
  assign _id2ex_io_Pc_NextD = pre_decoder_jump ? PCJumpD : _PC_nextD_T_2; // @[Mux.scala 101:16]
  assign _id2ex_io_BranchJump_JrD = {1'h0,__id2ex_io_BranchJump_JrD_T_2}; // @[Cat.scala 31:58]
  assign _if2id_clock = clk; // @[myCPU.scala 114:23]
  assign _if2id_reset = ~resetn; // @[myCPU.scala 114:41]
  assign _if2id_io_en = _cfu_io_StallD; // @[myCPU.scala 617:30]
  assign _if2id_io_clr = _cfu_io_FlushD; // @[myCPU.scala 618:30]
  assign _if2id_io_InstrF = {{32'd0}, __if2id_io_InstrF_T_5}; // @[myCPU.scala 621:27]
  assign _if2id_io_PCPlus4F = _if2id_io_PCF + 64'h4; // @[myCPU.scala 615:48]
  assign _if2id_io_PCF = fifo_with_bundle_io_read_out_0_pc; // @[myCPU.scala 602:36 603:26]
  assign _if2id_io_ExceptionTypeF = fifo_with_bundle_io_read_out_0_exception_type; // @[myCPU.scala 602:36 603:26]
  assign _mem22wb_clock = clk; // @[myCPU.scala 114:23]
  assign _mem22wb_reset = ~resetn; // @[myCPU.scala 114:41]
  assign _mem22wb_io_en = _cfu_io_StallW; // @[myCPU.scala 275:31]
  assign _mem22wb_io_clr = _cfu_io_FlushW; // @[myCPU.scala 276:31]
  assign _mem22wb_io_RegWriteM = _mem2mem2_io_RegWriteM; // @[myCPU.scala 278:38]
  assign _mem22wb_io_ResultM = _Forward_Lock1E_T_1 ? Mem_withRL_Data : ResultM2_Reg; // @[myCPU.scala 1105:25]
  assign _mem22wb_io_WriteRegM = _mem2mem2_io_WriteRegM; // @[myCPU.scala 280:38]
  assign _mem22wb_io_csrWriteM = _mem2mem2_io_csrWriteM; // @[myCPU.scala 282:38]
  assign _mem22wb_io_WritecsrAddrM = _mem2mem2_io_WritecsrAddrM; // @[myCPU.scala 283:38]
  assign _mem22wb_io_CsrWritedataM = _mem2mem2_io_CsrWritedataM; // @[myCPU.scala 1126:33]
  assign _mem22wb_io_PCM = _mem2mem2_io_PCM; // @[myCPU.scala 281:38]
  assign _mem22wb_io_ExceptionTypeM = _mem2mem2_io_ExceptionTypeM_Out; // @[myCPU.scala 1121:33]
  assign _mem22wb_io_BranchJump_JrM = _mem2mem2_io_BranchJump_JrM; // @[myCPU.scala 1125:33]
  assign _mem22wb_io_eBreakM = _mem2mem2_io_eBreakM; // @[myCPU.scala 1122:33]
  assign _mem22wb_io_Pc_NextM = _mem2mem2_io_Pc_NextM; // @[myCPU.scala 1123:33]
  assign _mem22wb_io_Mem_trace_budleM_pc = _mem2mem2_io_mem_trace_budleM_pc; // @[myCPU.scala 1130:37]
  assign _mem22wb_io_Mem_trace_budleM_data = __mem22wb_io_Mem_trace_budleM_data_T_2 |
    __mem22wb_io_Mem_trace_budleM_data_T_3; // @[Mux.scala 27:73]
  assign _mem22wb_io_Mem_trace_budleM_mem_fetch_type = _mem2mem2_io_mem_trace_budleM_mem_fetch_type; // @[myCPU.scala 1131:49]
  assign _mem22wb_io_Mem_trace_budleM_addr = _mem2mem2_io_mem_trace_budleM_addr; // @[myCPU.scala 1139:39]
  assign _mem22wb_io_Mem_trace_budleM_len = _mem2mem2_io_mem_trace_budleM_len; // @[myCPU.scala 1138:39]
  assign _mem22wb_io_Mem_trace_budleM_cache = _mem2mem2_io_mem_trace_budleM_cache; // @[myCPU.scala 1140:39]
  assign _addr_cal_io_d_vaddr = _id2ex_io_ImmE + RD1ForWardE; // @[myCPU.scala 1197:44]
  assign _muldiv_clock = clk; // @[myCPU.scala 114:23]
  assign _muldiv_reset = ~resetn; // @[myCPU.scala 114:41]
  assign _muldiv_io_en = ~ex_exception & ~__muldiv_io_en_T_23; // @[myCPU.scala 894:36]
  assign _muldiv_io_ctrl = _id2ex_io_muldiv_control; // @[myCPU.scala 901:21]
  assign _muldiv_io_in1 = _id2ex_io2_ALUSrcE_0 ? _id2ex_io2_PCE : RD1ForWardE; // @[myCPU.scala 876:20]
  assign _muldiv_io_in2 = _id2ex_io2_ALUSrcE_1 ? _id2ex_io_ImmE : RD2ForWardE; // @[myCPU.scala 883:20]
  assign _regfile_clock = clk; // @[myCPU.scala 114:23]
  assign _regfile_reset = ~resetn; // @[myCPU.scala 114:41]
  assign _regfile_io_A1 = _if2id_io_InstrD[19:15]; // @[myCPU.scala 769:29]
  assign _regfile_io_A2 = _if2id_io_InstrD[24:20]; // @[myCPU.scala 770:29]
  assign _regfile_io_WE3 = RegWriteW & _commit_difftest_data_ok_ok; // @[myCPU.scala 1169:41]
  assign _regfile_io_A3 = _mem22wb_io_WriteRegW; // @[myCPU.scala 1168:21]
  assign _regfile_io_WD3 = _mem22wb_io_ResultW; // @[myCPU.scala 1161:15 289:26]
  assign _mtrace_mod_reset = ~resetn; // @[myCPU.scala 227:29]
  assign _mtrace_mod_clock = clk; // @[myCPU.scala 226:26]
  assign _mtrace_mod_data = _mem22wb_io_Mem_trace_budleW_data; // @[myCPU.scala 236:29]
  assign _mtrace_mod_pc = _mem22wb_io_Mem_trace_budleW_pc; // @[myCPU.scala 228:26]
  assign _mtrace_mod_addr = _mem22wb_io_Mem_trace_budleW_addr; // @[myCPU.scala 234:29]
  assign _mtrace_mod_mem_req = _mem22wb_io_Mem_trace_budleW_mem_fetch_type != 2'h0; // @[myCPU.scala 229:75]
  assign _mtrace_mod_mem_write_read = _mem22wb_io_Mem_trace_budleW_mem_fetch_type[0]; // @[myCPU.scala 231:52]
  assign _mtrace_mod_mem_size = _mem22wb_io_Mem_trace_budleW_len; // @[myCPU.scala 235:29]
  assign _mtrace_mod_mem_cached = _mem22wb_io_Mem_trace_budleW_cache; // @[myCPU.scala 237:31]
  assign fifo_with_bundle_clock = clk; // @[myCPU.scala 114:23]
  assign fifo_with_bundle_reset = ~resetn; // @[myCPU.scala 114:41]
  assign fifo_with_bundle_io_read_en = {{1'd0}, _T_25}; // @[myCPU.scala 577:29]
  assign fifo_with_bundle_io_write_en = inst_write_en; // @[myCPU.scala 571:35]
  assign fifo_with_bundle_io_write_in_0_pc = stage_fec_2_pc_L_io_out_pc_value_out; // @[myCPU.scala 549:40 552:45]
  assign fifo_with_bundle_io_write_in_0_inst = inst_sram_rdata_L[31:0]; // @[myCPU.scala 551:60]
  assign fifo_with_bundle_io_write_in_0_pre_pc_target = branch_prediction_with_blockram_io_pre_target_L; // @[myCPU.scala 484:38 500:31]
  assign fifo_with_bundle_io_write_in_0_pre_lookup_data = branch_prediction_with_blockram_io_lookup_data_0; // @[myCPU.scala 487:40 489:29]
  assign fifo_with_bundle_io_write_in_0_pre_hashcode = stage_fec_2_hascode_0; // @[myCPU.scala 549:40 564:55]
  assign fifo_with_bundle_io_write_in_0_pre_pht = branch_prediction_with_blockram_io_out_L; // @[myCPU.scala 483:32 496:24]
  assign fifo_with_bundle_io_write_in_0_pre_bht = stage_fec_2_bht_0; // @[myCPU.scala 549:40 554:45]
  assign fifo_with_bundle_io_write_in_0_pre_lookup_value = branch_prediction_with_blockram_io_pht_lookup_value_out; // @[myCPU.scala 549:40 556:47]
  assign fifo_with_bundle_io_write_in_0_pre_decoder_branchD_flag = inst_sram_rdata_L[32]; // @[myCPU.scala 559:70]
  assign fifo_with_bundle_io_write_in_0_pre_decoder_jump = inst_sram_rdata_L[33]; // @[myCPU.scala 560:70]
  assign fifo_with_bundle_io_write_in_0_pre_decoder_branchdata = inst_sram_rdata_L[39:34]; // @[myCPU.scala 562:70]
  assign fifo_with_bundle_io_write_in_0_pre_decoder_jr = inst_buffer_write_bundle_pre_decoder_jr_opD == 7'h67 &
    inst_buffer_write_bundle_pre_decoder_jr_Funct3D == 3'h0; // @[macros.scala 497:30]
  assign fifo_with_bundle_io_write_in_0_true_branch_state = branch_prediction_with_blockram_io_pre_L & (
    stage_fec_2_inst_branch | stage_fec_2_inst_jump) & branch_prediction_with_blockram_io_btb_hit_0 &
    stage_fec_2_stall_reg & stage_fec_2_valid & ~_csr_io_exception; // @[myCPU.scala 511:187]
  assign fifo_with_bundle_io_point_write_en = _stage_fec_2_branch_answer_T_7 | _PCSrcD_T_1 & ((pre_decoder_jump |
    _PCSrcD_T_3) != id_true_branch_state | target_addr_error) & ~(ex_exception | mem_exception | mem2_exception |
    wb_exception); // @[myCPU.scala 732:60]
  assign fifo_with_bundle_io_point_flush = _csr_io_exception; // @[myCPU.scala 578:29]
  assign stage_fec_1_pc_L_clock = clk; // @[myCPU.scala 114:23]
  assign stage_fec_1_pc_L_reset = ~resetn; // @[myCPU.scala 114:41]
  assign stage_fec_1_pc_L_io_stall = stage2_stall; // @[myCPU.scala 444:31]
  assign stage_fec_1_pc_L_io_flush = _stage_fec_2_branch_answer_T_7 & ~stage2_stall; // @[myCPU.scala 402:54]
  assign stage_fec_1_pc_L_io_in_pc_value_in = _stage_fec_2_branch_answer_T_7 ? _csr_io_return_pc : _Pc_Next_T_3; // @[myCPU.scala 377:19]
  assign stage_fec_1_pc_M_clock = clk; // @[myCPU.scala 114:23]
  assign stage_fec_1_pc_M_reset = ~resetn; // @[myCPU.scala 114:41]
  assign stage_fec_1_pc_M_io_stall = stage2_stall; // @[myCPU.scala 445:31]
  assign stage_fec_1_pc_M_io_flush = _stage_fec_2_branch_answer_T_7 & ~stage2_stall; // @[myCPU.scala 402:54]
  assign stage_fec_1_pc_M_io_in_pc_value_in = _stage_fec_2_branch_answer_T_7 ? _csr_io_return_pc : _Pc_Next_T_3; // @[myCPU.scala 377:19]
  assign stage_fec_1_pc_R_clock = clk; // @[myCPU.scala 114:23]
  assign stage_fec_1_pc_R_reset = ~resetn; // @[myCPU.scala 114:41]
  assign stage_fec_1_pc_R_io_stall = stage2_stall; // @[myCPU.scala 446:31]
  assign stage_fec_1_pc_R_io_flush = _stage_fec_2_branch_answer_T_7 & ~stage2_stall; // @[myCPU.scala 402:54]
  assign stage_fec_1_pc_R_io_in_pc_value_in = _stage_fec_2_branch_answer_T_7 ? _csr_io_return_pc : _Pc_Next_T_3; // @[myCPU.scala 377:19]
  assign branch_prediction_with_blockram_clock = clk; // @[myCPU.scala 114:23]
  assign branch_prediction_with_blockram_reset = ~resetn; // @[myCPU.scala 114:41]
  assign branch_prediction_with_blockram_io_pc = stage_fec_1_pc_L_io_out_pc_value_out; // @[myCPU.scala 453:12]
  assign branch_prediction_with_blockram_io_write_pc = _mem22wb_io_PCW; // @[myCPU.scala 1186:17]
  assign branch_prediction_with_blockram_io_aw_pht_ways_addr = wb_bru_state_io_out_hashcode; // @[myCPU.scala 1185:25]
  assign branch_prediction_with_blockram_io_aw_pht_addr = wb_bru_state_io_out_lookup_data; // @[myCPU.scala 1183:20]
  assign branch_prediction_with_blockram_io_aw_bht_addr = _mem22wb_io_PCW[10:4]; // @[myCPU.scala 1182:38]
  assign branch_prediction_with_blockram_io_aw_target_addr = wb_bru_state_io_out_target_pc; // @[myCPU.scala 1184:23]
  assign branch_prediction_with_blockram_io_btb_write = branch_prediction_with_blockram_io_bht_write; // @[myCPU.scala 1181:18]
  assign branch_prediction_with_blockram_io_bht_write = _mem22wb_io_BranchJump_JrW[0]; // @[myCPU.scala 1179:47]
  assign branch_prediction_with_blockram_io_pht_write = branch_prediction_with_blockram_io_bht_write; // @[myCPU.scala 1180:18]
  assign branch_prediction_with_blockram_io_bht_in = wb_bru_state_io_out_bht; // @[myCPU.scala 1177:15]
  assign branch_prediction_with_blockram_io_pht_in = wb_bru_state_io_out_pht_lookup_value; // @[myCPU.scala 1178:15]
  assign branch_prediction_with_blockram_io_stage2_stall = stage2_stall & ~_pc_next_wait_T; // @[myCPU.scala 472:42]
  assign branch_prediction_with_blockram_io_stage2_flush = stage2_flush; // @[myCPU.scala 475:22]
  assign stage_fec_2_pc_L_clock = clk; // @[myCPU.scala 114:23]
  assign stage_fec_2_pc_L_reset = ~resetn; // @[myCPU.scala 114:41]
  assign stage_fec_2_pc_L_io_stall = stage2_stall & ~_pc_next_wait_T; // @[myCPU.scala 472:42]
  assign stage_fec_2_pc_L_io_flush = stage2_flush; // @[myCPU.scala 541:31]
  assign stage_fec_2_pc_L_io_in_pc_value_in = stage_fec_1_pc_L_io_out_pc_value_out; // @[myCPU.scala 532:40]
  assign stage_fec_2_pc_M_clock = clk; // @[myCPU.scala 114:23]
  assign stage_fec_2_pc_M_reset = ~resetn; // @[myCPU.scala 114:41]
  assign stage_fec_2_pc_M_io_stall = stage2_stall & ~_pc_next_wait_T; // @[myCPU.scala 472:42]
  assign stage_fec_2_pc_M_io_flush = stage2_flush; // @[myCPU.scala 542:31]
  assign stage_fec_2_pc_M_io_in_pc_value_in = stage_fec_1_pc_M_io_out_pc_value_out; // @[myCPU.scala 535:40]
  assign stage_fec_2_pc_R_clock = clk; // @[myCPU.scala 114:23]
  assign stage_fec_2_pc_R_reset = ~resetn; // @[myCPU.scala 114:41]
  assign stage_fec_2_pc_R_io_stall = stage2_stall & ~_pc_next_wait_T; // @[myCPU.scala 472:42]
  assign stage_fec_2_pc_R_io_flush = stage2_flush; // @[myCPU.scala 543:31]
  assign stage_fec_2_pc_R_io_in_pc_value_in = stage_fec_1_pc_R_io_out_pc_value_out; // @[myCPU.scala 538:40]
  assign id_bru_state_clock = clk; // @[myCPU.scala 114:23]
  assign id_bru_state_reset = ~resetn; // @[myCPU.scala 114:41]
  assign id_bru_state_io_stall = _cfu_io_StallD; // @[myCPU.scala 687:27]
  assign id_bru_state_io_flush = _cfu_io_FlushD; // @[myCPU.scala 686:27]
  assign id_bru_state_io_in_pht = fifo_with_bundle_io_read_out_0_pre_pht; // @[myCPU.scala 602:36 603:26]
  assign id_bru_state_io_in_bht = fifo_with_bundle_io_read_out_0_pre_bht; // @[myCPU.scala 602:36 603:26]
  assign id_bru_state_io_in_hashcode = fifo_with_bundle_io_read_out_0_pre_hashcode; // @[myCPU.scala 602:36 603:26]
  assign id_bru_state_io_in_target_pc = fifo_with_bundle_io_read_out_0_pre_pc_target; // @[myCPU.scala 602:36 603:26]
  assign id_bru_state_io_in_lookup_data = fifo_with_bundle_io_read_out_0_pre_lookup_data; // @[myCPU.scala 602:36 603:26]
  assign id_bru_state_io_in_pht_lookup_value = fifo_with_bundle_io_read_out_0_pre_lookup_value; // @[myCPU.scala 602:36 603:26]
  assign ex_bru_state_clock = clk; // @[myCPU.scala 114:23]
  assign ex_bru_state_reset = ~resetn; // @[myCPU.scala 114:41]
  assign ex_bru_state_io_stall = _cfu_io_StallE; // @[myCPU.scala 691:27]
  assign ex_bru_state_io_flush = _cfu_io_FlushE; // @[myCPU.scala 690:27]
  assign ex_bru_state_io_in_pht = id_bru_state_io_out_pht; // @[myCPU.scala 749:28]
  assign ex_bru_state_io_in_bht = id_bru_state_io_out_bht; // @[myCPU.scala 748:28]
  assign ex_bru_state_io_in_hashcode = id_bru_state_io_out_hashcode; // @[myCPU.scala 750:33]
  assign ex_bru_state_io_in_target_pc = pre_decoder_branchD_flag ? PCBranchD : _Pc_targetD_T_2; // @[Mux.scala 101:16]
  assign ex_bru_state_io_in_lookup_data = id_bru_state_io_out_lookup_data; // @[myCPU.scala 751:36]
  assign ex_bru_state_io_in_pht_lookup_value = id_bru_state_io_out_pht_lookup_value; // @[myCPU.scala 752:41]
  assign mem_bru_state_clock = clk; // @[myCPU.scala 114:23]
  assign mem_bru_state_reset = ~resetn; // @[myCPU.scala 114:41]
  assign mem_bru_state_io_stall = _cfu_io_StallM; // @[myCPU.scala 695:28]
  assign mem_bru_state_io_flush = _cfu_io_FlushM; // @[myCPU.scala 694:28]
  assign mem_bru_state_io_in_pht = 2'h2 == ex_bru_state_io_out_pht ? _pht_tobeE_T_3 : _pht_tobeE_T_7; // @[Mux.scala 81:58]
  assign mem_bru_state_io_in_bht = {ex_bru_state_io_out_bht[5:0],true_branch_stateE}; // @[Cat.scala 31:58]
  assign mem_bru_state_io_in_hashcode = ex_bru_state_io_out_hashcode; // @[myCPU.scala 706:26]
  assign mem_bru_state_io_in_target_pc = ex_bru_state_io_out_target_pc; // @[myCPU.scala 706:26]
  assign mem_bru_state_io_in_lookup_data = ex_bru_state_io_out_lookup_data; // @[myCPU.scala 706:26]
  assign mem_bru_state_io_in_pht_lookup_value = 2'h3 == ex_bru_state_io_out_lookup_data[1:0] ?
    _pht_lookup_value_tobeE_T_10 : _pht_lookup_value_tobeE_T_14; // @[Mux.scala 81:58]
  assign mem2_bru_state_clock = clk; // @[myCPU.scala 114:23]
  assign mem2_bru_state_reset = ~resetn; // @[myCPU.scala 114:41]
  assign mem2_bru_state_io_stall = _cfu_io_StallM2; // @[myCPU.scala 699:29]
  assign mem2_bru_state_io_flush = _cfu_io_FlushM2; // @[myCPU.scala 698:29]
  assign mem2_bru_state_io_in_pht = mem_bru_state_io_out_pht; // @[myCPU.scala 707:26]
  assign mem2_bru_state_io_in_bht = mem_bru_state_io_out_bht; // @[myCPU.scala 707:26]
  assign mem2_bru_state_io_in_hashcode = mem_bru_state_io_out_hashcode; // @[myCPU.scala 707:26]
  assign mem2_bru_state_io_in_target_pc = mem_bru_state_io_out_target_pc; // @[myCPU.scala 707:26]
  assign mem2_bru_state_io_in_lookup_data = mem_bru_state_io_out_lookup_data; // @[myCPU.scala 707:26]
  assign mem2_bru_state_io_in_pht_lookup_value = mem_bru_state_io_out_pht_lookup_value; // @[myCPU.scala 707:26]
  assign wb_bru_state_clock = clk; // @[myCPU.scala 114:23]
  assign wb_bru_state_reset = ~resetn; // @[myCPU.scala 114:41]
  assign wb_bru_state_io_stall = _cfu_io_StallW; // @[myCPU.scala 703:27]
  assign wb_bru_state_io_flush = _cfu_io_FlushW; // @[myCPU.scala 702:27]
  assign wb_bru_state_io_in_pht = mem2_bru_state_io_out_pht; // @[myCPU.scala 708:26]
  assign wb_bru_state_io_in_bht = mem2_bru_state_io_out_bht; // @[myCPU.scala 708:26]
  assign wb_bru_state_io_in_hashcode = mem2_bru_state_io_out_hashcode; // @[myCPU.scala 708:26]
  assign wb_bru_state_io_in_target_pc = mem2_bru_state_io_out_target_pc; // @[myCPU.scala 708:26]
  assign wb_bru_state_io_in_lookup_data = mem2_bru_state_io_out_lookup_data; // @[myCPU.scala 708:26]
  assign wb_bru_state_io_in_pht_lookup_value = mem2_bru_state_io_out_pht_lookup_value; // @[myCPU.scala 708:26]
  assign _commit_difftest_reset = ~resetn; // @[myCPU.scala 1150:34]
  assign _commit_difftest_clock = clk; // @[myCPU.scala 1149:31]
  assign _commit_difftest_gpr_wire = _regfile_io_reg_file_alL_out; // @[myCPU.scala 1151:34]
  assign _commit_difftest_pc = _mem22wb_io_PCW; // @[myCPU.scala 1153:40]
  assign _commit_difftest_debug_pc = wb_exception ? _csr_io_return_pc : _mem22wb_io_Pc_NextW; // @[myCPU.scala 1152:46]
  assign _commit_difftest_inst_commit = _PCW_Reg_T & pcw_reg != _mem22wb_io_PCW; // @[myCPU.scala 1159:64]
  assign _commit_difftest_cpu_ebreak_sign = _mem22wb_io_eBreakW; // @[myCPU.scala 1154:41]
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 606:36]
      pre_decoder_branchD_flag <= 1'h0;
    end else if (_cfu_io_FlushD) begin // @[myCPU.scala 606:66]
      pre_decoder_branchD_flag <= 1'h0;
    end else if (_PCSrcD_T_1) begin
      pre_decoder_branchD_flag <= inst_buffer_read_out_pre_decoder_branchD_flag;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 608:34]
      pre_decoder_branchdata <= 6'h0;
    end else if (_pre_decoder_branchD_flag_T) begin // @[myCPU.scala 608:64]
      pre_decoder_branchdata <= 6'h0;
    end else if (_PCSrcD_T_1) begin
      pre_decoder_branchdata <= inst_buffer_read_out_pre_decoder_branchdata;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 607:28]
      pre_decoder_jump <= 1'h0;
    end else if (_pre_decoder_branchD_flag_T) begin // @[myCPU.scala 607:58]
      pre_decoder_jump <= 1'h0;
    end else if (_PCSrcD_T_1) begin
      pre_decoder_jump <= inst_buffer_read_out_pre_decoder_jump;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 609:26]
      pre_decoder_jr <= 1'h0;
    end else if (_pre_decoder_branchD_flag_T) begin // @[myCPU.scala 609:56]
      pre_decoder_jr <= 1'h0;
    end else if (_PCSrcD_T_1) begin
      pre_decoder_jr <= inst_buffer_read_out_pre_decoder_jr;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 986:25]
      resultE2M_Reg <= 64'h0;
    end else if (_mem_exception_T) begin // @[myCPU.scala 986:55]
      resultE2M_Reg <= 64'h0;
    end else if (_mem_exception_T_1) begin
      resultE2M_Reg <= resultE;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 1037:24]
      ResultM2_Reg <= 64'h0;
    end else if (_mem2_exception_T) begin // @[myCPU.scala 1037:55]
      ResultM2_Reg <= 64'h0;
    end else if (_mem2_exception_T_1) begin
      ResultM2_Reg <= resultE2M_Reg;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 296:19]
      PCW_Reg <= 64'h0;
    end else if (_mem22wb_io_PCW != 64'h0) begin
      PCW_Reg <= _mem22wb_io_PCW;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 301:25]
      reg_pc <= 64'h0; // @[myCPU.scala 301:25]
    end else begin
      reg_pc <= _mem22wb_io_PCW; // @[myCPU.scala 302:12]
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 638:24]
      wb_exception <= 1'h0;
    end else if (_cfu_io_FlushW) begin // @[myCPU.scala 638:54]
      wb_exception <= 1'h0;
    end else if (_cfu_io_StallW) begin
      wb_exception <= _mem22wb_io_ExceptionTypeM != 32'h0;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 345:24]
      pc_next_wait <= 64'h0; // @[Mux.scala 101:{16,16} myCPU.scala 204:24 765:26 416:31]
    end else if (ready_to_branch | stage_fec_2_branch_answer) begin
      if (fifo_with_bundle_io_point_write_en) begin
        if (pre_decoder_jump) begin
          if (pre_decoder_jr) begin
            pc_next_wait <= _PCJumpD_T_58;
          end else begin
            pc_next_wait <= _PCJumpD_T_60;
          end
        end else if (_PCSrcD_T_3) begin
          pc_next_wait <= PCBranchD;
        end else begin
          pc_next_wait <= _if2id_io_PCPlus4D;
        end
      end else if (stage_fec_2_branch_answer) begin
        pc_next_wait <= stage_fec_2_pre_target_0;
      end else begin
        pc_next_wait <= _stage_fec_1_pc_next_T_1;
      end
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 472:42]
      stage_fec_2_stall_reg <= 1'h0;
    end else begin
      stage_fec_2_stall_reg <= stage2_stall & ~_pc_next_wait_T;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 480:29]
      stage_fec_2_valid <= 1'h0; // @[myCPU.scala 480:51]
    end else if (stage_fec_2_stall) begin
      if (fifo_with_bundle_io_point_write_en) begin
        stage_fec_2_valid <= 1'h0;
      end else begin
        stage_fec_2_valid <= stage_fec_1_valid;
      end
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 350:102]
      pc_req_wait <= 1'h0; // @[myCPU.scala 351:21]
    end else begin
      pc_req_wait <= ~inst_sram_en & _pc_next_wait_T & _stage_fec_2_branch_answer_T_8 | _GEN_0;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 360:28]
      exception_Pc_reg <= 64'h0;
    end else if (_stage_fec_2_branch_answer_T_7) begin
      exception_Pc_reg <= _csr_io_return_pc;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 365:58]
      returnPc_req_wait <= 1'h0; // @[myCPU.scala 366:27]
    end else begin
      returnPc_req_wait <= _T_4 & _stage_fec_2_branch_answer_T_7 | _GEN_2;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 462:29]
      stage_fec_1_valid <= 1'h0;
    end else begin
      stage_fec_1_valid <= stage2_stall | _stage_fec_1_valid_T_2;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 492:30]
      stage_fec_2_bht_0 <= 7'h0;
    end else if (stage2_flush) begin // @[myCPU.scala 492:51]
      stage_fec_2_bht_0 <= 7'h0;
    end else if (stage2_stall) begin
      stage_fec_2_bht_0 <= branch_prediction_with_blockram_io_bht_L;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 504:36]
      stage_fec_2_hascode_0 <= 4'h0;
    end else if (stage2_flush) begin // @[myCPU.scala 504:57]
      stage_fec_2_hascode_0 <= 4'h0;
    end else if (stage2_stall) begin
      stage_fec_2_hascode_0 <= _stage_fec_2_hascode_0_T_1;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 626:24]
      id_exception <= 1'h0;
    end else if (_pre_decoder_branchD_flag_T) begin // @[myCPU.scala 626:54]
      id_exception <= 1'h0;
    end else if (_PCSrcD_T_1) begin
      id_exception <= inst_buffer_read_out_pc[1:0] != 2'h0 | inst_buffer_read_out_exception_type != 2'h0;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 629:24]
      ex_exception <= 1'h0;
    end else if (_cfu_io_FlushE) begin // @[myCPU.scala 629:54]
      ex_exception <= 1'h0;
    end else if (_commit_cache_reg_T) begin
      ex_exception <= _id2ex_io_ExceptionTypeD != 32'h0;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 632:25]
      mem_exception <= 1'h0;
    end else if (_cfu_io_FlushM) begin // @[myCPU.scala 632:55]
      mem_exception <= 1'h0;
    end else if (_cfu_io_StallM) begin
      mem_exception <= _ex2mem_io_ExceptionTypeE != 32'h0;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 635:26]
      mem2_exception <= 1'h0;
    end else if (_cfu_io_FlushM2) begin // @[myCPU.scala 635:57]
      mem2_exception <= 1'h0;
    end else if (_cfu_io_StallM2) begin
      mem2_exception <= _mem2mem2_io_ExceptionTypeE != 32'h0;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 683:32]
      id_true_branch_state <= 1'h0;
    end else if (_pre_decoder_branchD_flag_T) begin // @[myCPU.scala 683:62]
      id_true_branch_state <= 1'h0;
    end else if (_PCSrcD_T_1) begin
      id_true_branch_state <= inst_buffer_read_out_true_branch_state;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 713:31]
      inst_tlb_exceptionE <= 1'h0;
    end else if (_ex_exception_T) begin // @[myCPU.scala 713:61]
      inst_tlb_exceptionE <= 1'h0;
    end else if (_commit_cache_reg_T) begin
      inst_tlb_exceptionE <= _if2id_io_ExceptionTypeD_Out != 2'h0;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 745:30]
      true_branch_stateE <= 1'h0;
    end else if (_ex_exception_T) begin // @[myCPU.scala 745:61]
      true_branch_stateE <= 1'h0;
    end else if (_commit_cache_reg_T) begin
      true_branch_stateE <= _T_31;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 793:25]
      int_instanceE_timer <= 1'h0;
    end else if (_ex_exception_T) begin // @[myCPU.scala 793:82]
      int_instanceE_timer <= 1'h0;
    end else if (_commit_cache_reg_T) begin
      int_instanceE_timer <= ext_int_timer;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 794:25]
      int_instanceM_timer <= 1'h0;
    end else if (_mem_exception_T) begin // @[myCPU.scala 794:82]
      int_instanceM_timer <= 1'h0;
    end else if (_mem_exception_T_1) begin
      int_instanceM_timer <= int_instanceE_timer;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 795:26]
      int_instanceM2_timer <= 1'h0;
    end else if (_mem2_exception_T) begin // @[myCPU.scala 795:82]
      int_instanceM2_timer <= 1'h0;
    end else if (_mem2_exception_T_1) begin
      int_instanceM2_timer <= int_instanceM_timer;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 796:25]
      int_instanceW_timer <= 1'h0;
    end else if (_wb_exception_T) begin // @[myCPU.scala 796:82]
      int_instanceW_timer <= 1'h0;
    end else if (_wb_exception_T_1) begin
      int_instanceW_timer <= int_instanceM2_timer;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 842:27]
      inst_tlb_exceptionM <= 1'h0;
    end else if (_mem_exception_T) begin // @[myCPU.scala 842:57]
      inst_tlb_exceptionM <= 1'h0;
    end else if (_mem_exception_T_1) begin
      inst_tlb_exceptionM <= inst_tlb_exceptionE;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 856:33]
      RD1ForWardE_r <= 64'h0; // @[myCPU.scala 846:34]
    end else if (!(_commit_cache_reg_T)) begin // @[myCPU.scala 860:88]
      if ((_cfu_io_Forward1E[0] | _cfu_io_Forward1E[1]) & ~Forward_Lock1E) begin // @[myCPU.scala 846:34]
        if (2'h3 == _cfu_io_Forward1E) begin
          RD1ForWardE_r <= ResultM2_Reg;
        end else if (2'h2 == _cfu_io_Forward1E) begin
          RD1ForWardE_r <= resultE2M_Reg;
        end else begin
          RD1ForWardE_r <= _RD1ForWardE_p_T_1;
        end
      end
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 856:33]
      RD2ForWardE_r <= 64'h0; // @[myCPU.scala 847:34]
    end else if (!(_commit_cache_reg_T)) begin // @[myCPU.scala 864:87]
      if ((_cfu_io_Forward2E[0] | _cfu_io_Forward2E[1]) & ~Forward_Lock2E) begin // @[myCPU.scala 847:34]
        if (2'h3 == _cfu_io_Forward2E) begin
          RD2ForWardE_r <= ResultM2_Reg;
        end else if (2'h2 == _cfu_io_Forward2E) begin
          RD2ForWardE_r <= resultE2M_Reg;
        end else begin
          RD2ForWardE_r <= _RD2ForWardE_p_T_1;
        end
      end
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 856:33]
      Forward_Lock1E <= 1'h0; // @[myCPU.scala 857:24]
    end else if (_commit_cache_reg_T) begin // @[myCPU.scala 860:88]
      Forward_Lock1E <= 1'h0; // @[myCPU.scala 861:28]
    end else if ((_cfu_io_Forward1E[0] | _cfu_io_Forward1E[1]) & ~Forward_Lock1E) begin // @[myCPU.scala 848:34]
      Forward_Lock1E <= ~(_ex2mem_io_MemToRegM | _mem2mem2_io_MemToRegM);
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 856:33]
      Forward_Lock2E <= 1'h0; // @[myCPU.scala 858:24]
    end else if (_commit_cache_reg_T) begin // @[myCPU.scala 864:87]
      Forward_Lock2E <= 1'h0; // @[myCPU.scala 865:28]
    end else if ((_cfu_io_Forward2E[0] | _cfu_io_Forward2E[1]) & ~Forward_Lock2E) begin // @[myCPU.scala 849:34]
      Forward_Lock2E <= _Forward_Lock1E_T_3;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 1085:33]
      tlb_exception_csr_writeM2 <= 1'h0;
    end else if (_mem2_exception_T) begin // @[myCPU.scala 1085:64]
      tlb_exception_csr_writeM2 <= 1'h0;
    end else if (_mem2_exception_T_1) begin
      tlb_exception_csr_writeM2 <= inst_tlb_exceptionM;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 1086:33]
      tlb_exception_co0_writeW <= 1'h0;
    end else if (_wb_exception_T) begin // @[myCPU.scala 1086:63]
      tlb_exception_co0_writeW <= 1'h0;
    end else if (_wb_exception_T_1) begin
      tlb_exception_co0_writeW <= tlb_exception_csr_writeM2;
    end
  end
  always @(posedge clk or posedge _T_2) begin
    if (_T_2) begin // @[myCPU.scala 1146:26]
      pcw_reg <= 64'h0; // @[myCPU.scala 1146:26]
    end else begin
      pcw_reg <= _mem22wb_io_PCW; // @[myCPU.scala 1156:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pre_decoder_branchD_flag = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  pre_decoder_branchdata = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  pre_decoder_jump = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  pre_decoder_jr = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  resultE2M_Reg = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  ResultM2_Reg = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  PCW_Reg = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  reg_pc = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  wb_exception = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  pc_next_wait = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  stage_fec_2_stall_reg = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  stage_fec_2_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  pc_req_wait = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  exception_Pc_reg = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  returnPc_req_wait = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  stage_fec_1_valid = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  stage_fec_2_bht_0 = _RAND_16[6:0];
  _RAND_17 = {1{`RANDOM}};
  stage_fec_2_hascode_0 = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  id_exception = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  ex_exception = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  mem_exception = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  mem2_exception = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  id_true_branch_state = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  inst_tlb_exceptionE = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  true_branch_stateE = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  int_instanceE_timer = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  int_instanceM_timer = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  int_instanceM2_timer = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  int_instanceW_timer = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  inst_tlb_exceptionM = _RAND_29[0:0];
  _RAND_30 = {2{`RANDOM}};
  RD1ForWardE_r = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  RD2ForWardE_r = _RAND_31[63:0];
  _RAND_32 = {1{`RANDOM}};
  Forward_Lock1E = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  Forward_Lock2E = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  tlb_exception_csr_writeM2 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  tlb_exception_co0_writeW = _RAND_35[0:0];
  _RAND_36 = {2{`RANDOM}};
  pcw_reg = _RAND_36[63:0];
`endif // RANDOMIZE_REG_INIT
  if (_T_2) begin
    pre_decoder_branchD_flag = 1'h0;
  end
  if (_T_2) begin
    pre_decoder_branchdata = 6'h0;
  end
  if (_T_2) begin
    pre_decoder_jump = 1'h0;
  end
  if (_T_2) begin
    pre_decoder_jr = 1'h0;
  end
  if (_T_2) begin
    resultE2M_Reg = 64'h0;
  end
  if (_T_2) begin
    ResultM2_Reg = 64'h0;
  end
  if (_T_2) begin
    PCW_Reg = 64'h0;
  end
  if (_T_2) begin
    reg_pc = 64'h0;
  end
  if (_T_2) begin
    wb_exception = 1'h0;
  end
  if (_T_2) begin
    pc_next_wait = 64'h0;
  end
  if (_T_2) begin
    stage_fec_2_stall_reg = 1'h0;
  end
  if (_T_2) begin
    stage_fec_2_valid = 1'h0;
  end
  if (_T_2) begin
    pc_req_wait = 1'h0;
  end
  if (_T_2) begin
    exception_Pc_reg = 64'h0;
  end
  if (_T_2) begin
    returnPc_req_wait = 1'h0;
  end
  if (_T_2) begin
    stage_fec_1_valid = 1'h0;
  end
  if (_T_2) begin
    stage_fec_2_bht_0 = 7'h0;
  end
  if (_T_2) begin
    stage_fec_2_hascode_0 = 4'h0;
  end
  if (_T_2) begin
    id_exception = 1'h0;
  end
  if (_T_2) begin
    ex_exception = 1'h0;
  end
  if (_T_2) begin
    mem_exception = 1'h0;
  end
  if (_T_2) begin
    mem2_exception = 1'h0;
  end
  if (_T_2) begin
    id_true_branch_state = 1'h0;
  end
  if (_T_2) begin
    inst_tlb_exceptionE = 1'h0;
  end
  if (_T_2) begin
    true_branch_stateE = 1'h0;
  end
  if (_T_2) begin
    int_instanceE_timer = 1'h0;
  end
  if (_T_2) begin
    int_instanceM_timer = 1'h0;
  end
  if (_T_2) begin
    int_instanceM2_timer = 1'h0;
  end
  if (_T_2) begin
    int_instanceW_timer = 1'h0;
  end
  if (_T_2) begin
    inst_tlb_exceptionM = 1'h0;
  end
  if (_T_2) begin
    RD1ForWardE_r = 64'h0;
  end
  if (_T_2) begin
    RD2ForWardE_r = 64'h0;
  end
  if (_T_2) begin
    Forward_Lock1E = 1'h0;
  end
  if (_T_2) begin
    Forward_Lock2E = 1'h0;
  end
  if (_T_2) begin
    tlb_exception_csr_writeM2 = 1'h0;
  end
  if (_T_2) begin
    tlb_exception_co0_writeW = 1'h0;
  end
  if (_T_2) begin
    pcw_reg = 64'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module icache_tag(
  input         clock,
  input         reset,
  input         io_wen,
  input  [20:0] io_wdata,
  input  [63:0] io_addr,
  output        io_hit,
  output        io_valid,
  input         io_tag_all_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
`endif // RANDOMIZE_REG_INIT
  reg [21:0] tag_regs_0; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_1; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_2; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_3; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_4; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_5; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_6; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_7; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_8; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_9; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_10; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_11; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_12; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_13; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_14; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_15; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_16; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_17; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_18; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_19; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_20; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_21; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_22; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_23; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_24; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_25; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_26; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_27; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_28; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_29; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_30; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_31; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_32; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_33; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_34; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_35; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_36; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_37; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_38; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_39; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_40; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_41; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_42; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_43; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_44; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_45; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_46; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_47; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_48; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_49; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_50; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_51; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_52; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_53; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_54; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_55; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_56; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_57; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_58; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_59; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_60; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_61; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_62; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_63; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_64; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_65; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_66; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_67; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_68; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_69; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_70; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_71; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_72; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_73; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_74; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_75; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_76; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_77; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_78; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_79; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_80; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_81; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_82; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_83; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_84; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_85; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_86; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_87; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_88; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_89; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_90; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_91; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_92; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_93; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_94; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_95; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_96; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_97; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_98; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_99; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_100; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_101; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_102; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_103; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_104; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_105; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_106; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_107; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_108; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_109; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_110; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_111; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_112; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_113; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_114; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_115; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_116; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_117; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_118; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_119; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_120; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_121; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_122; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_123; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_124; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_125; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_126; // @[icache_tag.scala 21:27]
  reg [21:0] tag_regs_127; // @[icache_tag.scala 21:27]
  reg [7:0] tag_asid_regs_0; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_1; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_2; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_3; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_4; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_5; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_6; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_7; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_8; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_9; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_10; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_11; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_12; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_13; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_14; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_15; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_16; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_17; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_18; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_19; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_20; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_21; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_22; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_23; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_24; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_25; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_26; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_27; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_28; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_29; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_30; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_31; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_32; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_33; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_34; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_35; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_36; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_37; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_38; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_39; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_40; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_41; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_42; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_43; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_44; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_45; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_46; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_47; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_48; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_49; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_50; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_51; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_52; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_53; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_54; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_55; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_56; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_57; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_58; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_59; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_60; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_61; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_62; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_63; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_64; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_65; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_66; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_67; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_68; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_69; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_70; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_71; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_72; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_73; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_74; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_75; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_76; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_77; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_78; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_79; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_80; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_81; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_82; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_83; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_84; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_85; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_86; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_87; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_88; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_89; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_90; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_91; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_92; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_93; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_94; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_95; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_96; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_97; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_98; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_99; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_100; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_101; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_102; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_103; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_104; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_105; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_106; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_107; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_108; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_109; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_110; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_111; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_112; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_113; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_114; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_115; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_116; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_117; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_118; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_119; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_120; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_121; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_122; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_123; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_124; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_125; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_126; // @[icache_tag.scala 22:32]
  reg [7:0] tag_asid_regs_127; // @[icache_tag.scala 22:32]
  wire  _valid_to_be_T_5 = io_wen & io_addr[10:4] == 7'h0; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_8 = io_wen & io_addr[10:4] == 7'h0 ? io_wdata[20] : tag_regs_0[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be = io_tag_all_flush ? 1'h0 : _valid_to_be_T_8; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be = _valid_to_be_T_5 ? io_wdata[19:0] : tag_regs_0[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_0_T = {valid_to_be,tag_to_be}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_14 = io_wen & io_addr[10:4] == 7'h1; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_17 = io_wen & io_addr[10:4] == 7'h1 ? io_wdata[20] : tag_regs_1[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_1 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_17; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_1 = _valid_to_be_T_14 ? io_wdata[19:0] : tag_regs_1[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_1_T = {valid_to_be_1,tag_to_be_1}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_23 = io_wen & io_addr[10:4] == 7'h2; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_26 = io_wen & io_addr[10:4] == 7'h2 ? io_wdata[20] : tag_regs_2[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_2 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_26; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_2 = _valid_to_be_T_23 ? io_wdata[19:0] : tag_regs_2[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_2_T = {valid_to_be_2,tag_to_be_2}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_32 = io_wen & io_addr[10:4] == 7'h3; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_35 = io_wen & io_addr[10:4] == 7'h3 ? io_wdata[20] : tag_regs_3[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_3 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_35; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_3 = _valid_to_be_T_32 ? io_wdata[19:0] : tag_regs_3[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_3_T = {valid_to_be_3,tag_to_be_3}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_41 = io_wen & io_addr[10:4] == 7'h4; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_44 = io_wen & io_addr[10:4] == 7'h4 ? io_wdata[20] : tag_regs_4[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_4 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_44; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_4 = _valid_to_be_T_41 ? io_wdata[19:0] : tag_regs_4[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_4_T = {valid_to_be_4,tag_to_be_4}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_50 = io_wen & io_addr[10:4] == 7'h5; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_53 = io_wen & io_addr[10:4] == 7'h5 ? io_wdata[20] : tag_regs_5[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_5 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_53; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_5 = _valid_to_be_T_50 ? io_wdata[19:0] : tag_regs_5[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_5_T = {valid_to_be_5,tag_to_be_5}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_59 = io_wen & io_addr[10:4] == 7'h6; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_62 = io_wen & io_addr[10:4] == 7'h6 ? io_wdata[20] : tag_regs_6[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_6 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_62; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_6 = _valid_to_be_T_59 ? io_wdata[19:0] : tag_regs_6[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_6_T = {valid_to_be_6,tag_to_be_6}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_68 = io_wen & io_addr[10:4] == 7'h7; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_71 = io_wen & io_addr[10:4] == 7'h7 ? io_wdata[20] : tag_regs_7[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_7 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_71; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_7 = _valid_to_be_T_68 ? io_wdata[19:0] : tag_regs_7[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_7_T = {valid_to_be_7,tag_to_be_7}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_77 = io_wen & io_addr[10:4] == 7'h8; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_80 = io_wen & io_addr[10:4] == 7'h8 ? io_wdata[20] : tag_regs_8[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_8 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_80; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_8 = _valid_to_be_T_77 ? io_wdata[19:0] : tag_regs_8[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_8_T = {valid_to_be_8,tag_to_be_8}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_86 = io_wen & io_addr[10:4] == 7'h9; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_89 = io_wen & io_addr[10:4] == 7'h9 ? io_wdata[20] : tag_regs_9[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_9 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_89; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_9 = _valid_to_be_T_86 ? io_wdata[19:0] : tag_regs_9[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_9_T = {valid_to_be_9,tag_to_be_9}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_95 = io_wen & io_addr[10:4] == 7'ha; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_98 = io_wen & io_addr[10:4] == 7'ha ? io_wdata[20] : tag_regs_10[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_10 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_98; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_10 = _valid_to_be_T_95 ? io_wdata[19:0] : tag_regs_10[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_10_T = {valid_to_be_10,tag_to_be_10}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_104 = io_wen & io_addr[10:4] == 7'hb; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_107 = io_wen & io_addr[10:4] == 7'hb ? io_wdata[20] : tag_regs_11[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_11 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_107; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_11 = _valid_to_be_T_104 ? io_wdata[19:0] : tag_regs_11[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_11_T = {valid_to_be_11,tag_to_be_11}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_113 = io_wen & io_addr[10:4] == 7'hc; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_116 = io_wen & io_addr[10:4] == 7'hc ? io_wdata[20] : tag_regs_12[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_12 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_116; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_12 = _valid_to_be_T_113 ? io_wdata[19:0] : tag_regs_12[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_12_T = {valid_to_be_12,tag_to_be_12}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_122 = io_wen & io_addr[10:4] == 7'hd; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_125 = io_wen & io_addr[10:4] == 7'hd ? io_wdata[20] : tag_regs_13[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_13 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_125; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_13 = _valid_to_be_T_122 ? io_wdata[19:0] : tag_regs_13[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_13_T = {valid_to_be_13,tag_to_be_13}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_131 = io_wen & io_addr[10:4] == 7'he; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_134 = io_wen & io_addr[10:4] == 7'he ? io_wdata[20] : tag_regs_14[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_14 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_134; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_14 = _valid_to_be_T_131 ? io_wdata[19:0] : tag_regs_14[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_14_T = {valid_to_be_14,tag_to_be_14}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_140 = io_wen & io_addr[10:4] == 7'hf; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_143 = io_wen & io_addr[10:4] == 7'hf ? io_wdata[20] : tag_regs_15[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_15 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_143; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_15 = _valid_to_be_T_140 ? io_wdata[19:0] : tag_regs_15[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_15_T = {valid_to_be_15,tag_to_be_15}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_149 = io_wen & io_addr[10:4] == 7'h10; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_152 = io_wen & io_addr[10:4] == 7'h10 ? io_wdata[20] : tag_regs_16[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_16 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_152; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_16 = _valid_to_be_T_149 ? io_wdata[19:0] : tag_regs_16[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_16_T = {valid_to_be_16,tag_to_be_16}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_158 = io_wen & io_addr[10:4] == 7'h11; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_161 = io_wen & io_addr[10:4] == 7'h11 ? io_wdata[20] : tag_regs_17[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_17 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_161; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_17 = _valid_to_be_T_158 ? io_wdata[19:0] : tag_regs_17[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_17_T = {valid_to_be_17,tag_to_be_17}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_167 = io_wen & io_addr[10:4] == 7'h12; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_170 = io_wen & io_addr[10:4] == 7'h12 ? io_wdata[20] : tag_regs_18[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_18 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_170; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_18 = _valid_to_be_T_167 ? io_wdata[19:0] : tag_regs_18[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_18_T = {valid_to_be_18,tag_to_be_18}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_176 = io_wen & io_addr[10:4] == 7'h13; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_179 = io_wen & io_addr[10:4] == 7'h13 ? io_wdata[20] : tag_regs_19[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_19 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_179; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_19 = _valid_to_be_T_176 ? io_wdata[19:0] : tag_regs_19[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_19_T = {valid_to_be_19,tag_to_be_19}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_185 = io_wen & io_addr[10:4] == 7'h14; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_188 = io_wen & io_addr[10:4] == 7'h14 ? io_wdata[20] : tag_regs_20[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_20 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_188; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_20 = _valid_to_be_T_185 ? io_wdata[19:0] : tag_regs_20[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_20_T = {valid_to_be_20,tag_to_be_20}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_194 = io_wen & io_addr[10:4] == 7'h15; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_197 = io_wen & io_addr[10:4] == 7'h15 ? io_wdata[20] : tag_regs_21[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_21 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_197; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_21 = _valid_to_be_T_194 ? io_wdata[19:0] : tag_regs_21[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_21_T = {valid_to_be_21,tag_to_be_21}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_203 = io_wen & io_addr[10:4] == 7'h16; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_206 = io_wen & io_addr[10:4] == 7'h16 ? io_wdata[20] : tag_regs_22[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_22 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_206; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_22 = _valid_to_be_T_203 ? io_wdata[19:0] : tag_regs_22[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_22_T = {valid_to_be_22,tag_to_be_22}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_212 = io_wen & io_addr[10:4] == 7'h17; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_215 = io_wen & io_addr[10:4] == 7'h17 ? io_wdata[20] : tag_regs_23[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_23 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_215; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_23 = _valid_to_be_T_212 ? io_wdata[19:0] : tag_regs_23[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_23_T = {valid_to_be_23,tag_to_be_23}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_221 = io_wen & io_addr[10:4] == 7'h18; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_224 = io_wen & io_addr[10:4] == 7'h18 ? io_wdata[20] : tag_regs_24[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_24 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_224; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_24 = _valid_to_be_T_221 ? io_wdata[19:0] : tag_regs_24[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_24_T = {valid_to_be_24,tag_to_be_24}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_230 = io_wen & io_addr[10:4] == 7'h19; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_233 = io_wen & io_addr[10:4] == 7'h19 ? io_wdata[20] : tag_regs_25[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_25 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_233; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_25 = _valid_to_be_T_230 ? io_wdata[19:0] : tag_regs_25[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_25_T = {valid_to_be_25,tag_to_be_25}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_239 = io_wen & io_addr[10:4] == 7'h1a; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_242 = io_wen & io_addr[10:4] == 7'h1a ? io_wdata[20] : tag_regs_26[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_26 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_242; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_26 = _valid_to_be_T_239 ? io_wdata[19:0] : tag_regs_26[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_26_T = {valid_to_be_26,tag_to_be_26}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_248 = io_wen & io_addr[10:4] == 7'h1b; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_251 = io_wen & io_addr[10:4] == 7'h1b ? io_wdata[20] : tag_regs_27[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_27 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_251; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_27 = _valid_to_be_T_248 ? io_wdata[19:0] : tag_regs_27[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_27_T = {valid_to_be_27,tag_to_be_27}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_257 = io_wen & io_addr[10:4] == 7'h1c; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_260 = io_wen & io_addr[10:4] == 7'h1c ? io_wdata[20] : tag_regs_28[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_28 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_260; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_28 = _valid_to_be_T_257 ? io_wdata[19:0] : tag_regs_28[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_28_T = {valid_to_be_28,tag_to_be_28}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_266 = io_wen & io_addr[10:4] == 7'h1d; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_269 = io_wen & io_addr[10:4] == 7'h1d ? io_wdata[20] : tag_regs_29[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_29 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_269; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_29 = _valid_to_be_T_266 ? io_wdata[19:0] : tag_regs_29[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_29_T = {valid_to_be_29,tag_to_be_29}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_275 = io_wen & io_addr[10:4] == 7'h1e; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_278 = io_wen & io_addr[10:4] == 7'h1e ? io_wdata[20] : tag_regs_30[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_30 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_278; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_30 = _valid_to_be_T_275 ? io_wdata[19:0] : tag_regs_30[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_30_T = {valid_to_be_30,tag_to_be_30}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_284 = io_wen & io_addr[10:4] == 7'h1f; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_287 = io_wen & io_addr[10:4] == 7'h1f ? io_wdata[20] : tag_regs_31[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_31 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_287; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_31 = _valid_to_be_T_284 ? io_wdata[19:0] : tag_regs_31[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_31_T = {valid_to_be_31,tag_to_be_31}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_293 = io_wen & io_addr[10:4] == 7'h20; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_296 = io_wen & io_addr[10:4] == 7'h20 ? io_wdata[20] : tag_regs_32[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_32 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_296; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_32 = _valid_to_be_T_293 ? io_wdata[19:0] : tag_regs_32[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_32_T = {valid_to_be_32,tag_to_be_32}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_302 = io_wen & io_addr[10:4] == 7'h21; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_305 = io_wen & io_addr[10:4] == 7'h21 ? io_wdata[20] : tag_regs_33[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_33 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_305; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_33 = _valid_to_be_T_302 ? io_wdata[19:0] : tag_regs_33[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_33_T = {valid_to_be_33,tag_to_be_33}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_311 = io_wen & io_addr[10:4] == 7'h22; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_314 = io_wen & io_addr[10:4] == 7'h22 ? io_wdata[20] : tag_regs_34[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_34 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_314; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_34 = _valid_to_be_T_311 ? io_wdata[19:0] : tag_regs_34[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_34_T = {valid_to_be_34,tag_to_be_34}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_320 = io_wen & io_addr[10:4] == 7'h23; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_323 = io_wen & io_addr[10:4] == 7'h23 ? io_wdata[20] : tag_regs_35[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_35 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_323; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_35 = _valid_to_be_T_320 ? io_wdata[19:0] : tag_regs_35[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_35_T = {valid_to_be_35,tag_to_be_35}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_329 = io_wen & io_addr[10:4] == 7'h24; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_332 = io_wen & io_addr[10:4] == 7'h24 ? io_wdata[20] : tag_regs_36[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_36 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_332; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_36 = _valid_to_be_T_329 ? io_wdata[19:0] : tag_regs_36[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_36_T = {valid_to_be_36,tag_to_be_36}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_338 = io_wen & io_addr[10:4] == 7'h25; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_341 = io_wen & io_addr[10:4] == 7'h25 ? io_wdata[20] : tag_regs_37[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_37 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_341; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_37 = _valid_to_be_T_338 ? io_wdata[19:0] : tag_regs_37[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_37_T = {valid_to_be_37,tag_to_be_37}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_347 = io_wen & io_addr[10:4] == 7'h26; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_350 = io_wen & io_addr[10:4] == 7'h26 ? io_wdata[20] : tag_regs_38[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_38 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_350; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_38 = _valid_to_be_T_347 ? io_wdata[19:0] : tag_regs_38[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_38_T = {valid_to_be_38,tag_to_be_38}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_356 = io_wen & io_addr[10:4] == 7'h27; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_359 = io_wen & io_addr[10:4] == 7'h27 ? io_wdata[20] : tag_regs_39[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_39 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_359; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_39 = _valid_to_be_T_356 ? io_wdata[19:0] : tag_regs_39[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_39_T = {valid_to_be_39,tag_to_be_39}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_365 = io_wen & io_addr[10:4] == 7'h28; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_368 = io_wen & io_addr[10:4] == 7'h28 ? io_wdata[20] : tag_regs_40[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_40 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_368; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_40 = _valid_to_be_T_365 ? io_wdata[19:0] : tag_regs_40[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_40_T = {valid_to_be_40,tag_to_be_40}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_374 = io_wen & io_addr[10:4] == 7'h29; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_377 = io_wen & io_addr[10:4] == 7'h29 ? io_wdata[20] : tag_regs_41[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_41 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_377; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_41 = _valid_to_be_T_374 ? io_wdata[19:0] : tag_regs_41[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_41_T = {valid_to_be_41,tag_to_be_41}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_383 = io_wen & io_addr[10:4] == 7'h2a; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_386 = io_wen & io_addr[10:4] == 7'h2a ? io_wdata[20] : tag_regs_42[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_42 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_386; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_42 = _valid_to_be_T_383 ? io_wdata[19:0] : tag_regs_42[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_42_T = {valid_to_be_42,tag_to_be_42}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_392 = io_wen & io_addr[10:4] == 7'h2b; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_395 = io_wen & io_addr[10:4] == 7'h2b ? io_wdata[20] : tag_regs_43[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_43 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_395; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_43 = _valid_to_be_T_392 ? io_wdata[19:0] : tag_regs_43[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_43_T = {valid_to_be_43,tag_to_be_43}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_401 = io_wen & io_addr[10:4] == 7'h2c; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_404 = io_wen & io_addr[10:4] == 7'h2c ? io_wdata[20] : tag_regs_44[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_44 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_404; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_44 = _valid_to_be_T_401 ? io_wdata[19:0] : tag_regs_44[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_44_T = {valid_to_be_44,tag_to_be_44}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_410 = io_wen & io_addr[10:4] == 7'h2d; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_413 = io_wen & io_addr[10:4] == 7'h2d ? io_wdata[20] : tag_regs_45[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_45 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_413; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_45 = _valid_to_be_T_410 ? io_wdata[19:0] : tag_regs_45[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_45_T = {valid_to_be_45,tag_to_be_45}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_419 = io_wen & io_addr[10:4] == 7'h2e; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_422 = io_wen & io_addr[10:4] == 7'h2e ? io_wdata[20] : tag_regs_46[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_46 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_422; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_46 = _valid_to_be_T_419 ? io_wdata[19:0] : tag_regs_46[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_46_T = {valid_to_be_46,tag_to_be_46}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_428 = io_wen & io_addr[10:4] == 7'h2f; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_431 = io_wen & io_addr[10:4] == 7'h2f ? io_wdata[20] : tag_regs_47[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_47 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_431; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_47 = _valid_to_be_T_428 ? io_wdata[19:0] : tag_regs_47[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_47_T = {valid_to_be_47,tag_to_be_47}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_437 = io_wen & io_addr[10:4] == 7'h30; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_440 = io_wen & io_addr[10:4] == 7'h30 ? io_wdata[20] : tag_regs_48[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_48 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_440; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_48 = _valid_to_be_T_437 ? io_wdata[19:0] : tag_regs_48[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_48_T = {valid_to_be_48,tag_to_be_48}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_446 = io_wen & io_addr[10:4] == 7'h31; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_449 = io_wen & io_addr[10:4] == 7'h31 ? io_wdata[20] : tag_regs_49[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_49 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_449; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_49 = _valid_to_be_T_446 ? io_wdata[19:0] : tag_regs_49[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_49_T = {valid_to_be_49,tag_to_be_49}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_455 = io_wen & io_addr[10:4] == 7'h32; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_458 = io_wen & io_addr[10:4] == 7'h32 ? io_wdata[20] : tag_regs_50[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_50 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_458; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_50 = _valid_to_be_T_455 ? io_wdata[19:0] : tag_regs_50[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_50_T = {valid_to_be_50,tag_to_be_50}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_464 = io_wen & io_addr[10:4] == 7'h33; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_467 = io_wen & io_addr[10:4] == 7'h33 ? io_wdata[20] : tag_regs_51[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_51 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_467; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_51 = _valid_to_be_T_464 ? io_wdata[19:0] : tag_regs_51[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_51_T = {valid_to_be_51,tag_to_be_51}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_473 = io_wen & io_addr[10:4] == 7'h34; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_476 = io_wen & io_addr[10:4] == 7'h34 ? io_wdata[20] : tag_regs_52[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_52 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_476; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_52 = _valid_to_be_T_473 ? io_wdata[19:0] : tag_regs_52[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_52_T = {valid_to_be_52,tag_to_be_52}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_482 = io_wen & io_addr[10:4] == 7'h35; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_485 = io_wen & io_addr[10:4] == 7'h35 ? io_wdata[20] : tag_regs_53[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_53 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_485; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_53 = _valid_to_be_T_482 ? io_wdata[19:0] : tag_regs_53[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_53_T = {valid_to_be_53,tag_to_be_53}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_491 = io_wen & io_addr[10:4] == 7'h36; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_494 = io_wen & io_addr[10:4] == 7'h36 ? io_wdata[20] : tag_regs_54[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_54 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_494; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_54 = _valid_to_be_T_491 ? io_wdata[19:0] : tag_regs_54[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_54_T = {valid_to_be_54,tag_to_be_54}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_500 = io_wen & io_addr[10:4] == 7'h37; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_503 = io_wen & io_addr[10:4] == 7'h37 ? io_wdata[20] : tag_regs_55[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_55 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_503; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_55 = _valid_to_be_T_500 ? io_wdata[19:0] : tag_regs_55[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_55_T = {valid_to_be_55,tag_to_be_55}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_509 = io_wen & io_addr[10:4] == 7'h38; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_512 = io_wen & io_addr[10:4] == 7'h38 ? io_wdata[20] : tag_regs_56[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_56 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_512; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_56 = _valid_to_be_T_509 ? io_wdata[19:0] : tag_regs_56[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_56_T = {valid_to_be_56,tag_to_be_56}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_518 = io_wen & io_addr[10:4] == 7'h39; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_521 = io_wen & io_addr[10:4] == 7'h39 ? io_wdata[20] : tag_regs_57[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_57 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_521; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_57 = _valid_to_be_T_518 ? io_wdata[19:0] : tag_regs_57[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_57_T = {valid_to_be_57,tag_to_be_57}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_527 = io_wen & io_addr[10:4] == 7'h3a; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_530 = io_wen & io_addr[10:4] == 7'h3a ? io_wdata[20] : tag_regs_58[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_58 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_530; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_58 = _valid_to_be_T_527 ? io_wdata[19:0] : tag_regs_58[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_58_T = {valid_to_be_58,tag_to_be_58}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_536 = io_wen & io_addr[10:4] == 7'h3b; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_539 = io_wen & io_addr[10:4] == 7'h3b ? io_wdata[20] : tag_regs_59[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_59 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_539; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_59 = _valid_to_be_T_536 ? io_wdata[19:0] : tag_regs_59[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_59_T = {valid_to_be_59,tag_to_be_59}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_545 = io_wen & io_addr[10:4] == 7'h3c; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_548 = io_wen & io_addr[10:4] == 7'h3c ? io_wdata[20] : tag_regs_60[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_60 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_548; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_60 = _valid_to_be_T_545 ? io_wdata[19:0] : tag_regs_60[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_60_T = {valid_to_be_60,tag_to_be_60}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_554 = io_wen & io_addr[10:4] == 7'h3d; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_557 = io_wen & io_addr[10:4] == 7'h3d ? io_wdata[20] : tag_regs_61[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_61 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_557; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_61 = _valid_to_be_T_554 ? io_wdata[19:0] : tag_regs_61[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_61_T = {valid_to_be_61,tag_to_be_61}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_563 = io_wen & io_addr[10:4] == 7'h3e; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_566 = io_wen & io_addr[10:4] == 7'h3e ? io_wdata[20] : tag_regs_62[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_62 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_566; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_62 = _valid_to_be_T_563 ? io_wdata[19:0] : tag_regs_62[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_62_T = {valid_to_be_62,tag_to_be_62}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_572 = io_wen & io_addr[10:4] == 7'h3f; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_575 = io_wen & io_addr[10:4] == 7'h3f ? io_wdata[20] : tag_regs_63[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_63 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_575; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_63 = _valid_to_be_T_572 ? io_wdata[19:0] : tag_regs_63[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_63_T = {valid_to_be_63,tag_to_be_63}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_581 = io_wen & io_addr[10:4] == 7'h40; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_584 = io_wen & io_addr[10:4] == 7'h40 ? io_wdata[20] : tag_regs_64[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_64 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_584; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_64 = _valid_to_be_T_581 ? io_wdata[19:0] : tag_regs_64[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_64_T = {valid_to_be_64,tag_to_be_64}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_590 = io_wen & io_addr[10:4] == 7'h41; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_593 = io_wen & io_addr[10:4] == 7'h41 ? io_wdata[20] : tag_regs_65[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_65 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_593; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_65 = _valid_to_be_T_590 ? io_wdata[19:0] : tag_regs_65[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_65_T = {valid_to_be_65,tag_to_be_65}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_599 = io_wen & io_addr[10:4] == 7'h42; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_602 = io_wen & io_addr[10:4] == 7'h42 ? io_wdata[20] : tag_regs_66[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_66 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_602; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_66 = _valid_to_be_T_599 ? io_wdata[19:0] : tag_regs_66[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_66_T = {valid_to_be_66,tag_to_be_66}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_608 = io_wen & io_addr[10:4] == 7'h43; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_611 = io_wen & io_addr[10:4] == 7'h43 ? io_wdata[20] : tag_regs_67[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_67 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_611; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_67 = _valid_to_be_T_608 ? io_wdata[19:0] : tag_regs_67[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_67_T = {valid_to_be_67,tag_to_be_67}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_617 = io_wen & io_addr[10:4] == 7'h44; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_620 = io_wen & io_addr[10:4] == 7'h44 ? io_wdata[20] : tag_regs_68[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_68 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_620; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_68 = _valid_to_be_T_617 ? io_wdata[19:0] : tag_regs_68[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_68_T = {valid_to_be_68,tag_to_be_68}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_626 = io_wen & io_addr[10:4] == 7'h45; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_629 = io_wen & io_addr[10:4] == 7'h45 ? io_wdata[20] : tag_regs_69[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_69 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_629; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_69 = _valid_to_be_T_626 ? io_wdata[19:0] : tag_regs_69[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_69_T = {valid_to_be_69,tag_to_be_69}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_635 = io_wen & io_addr[10:4] == 7'h46; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_638 = io_wen & io_addr[10:4] == 7'h46 ? io_wdata[20] : tag_regs_70[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_70 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_638; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_70 = _valid_to_be_T_635 ? io_wdata[19:0] : tag_regs_70[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_70_T = {valid_to_be_70,tag_to_be_70}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_644 = io_wen & io_addr[10:4] == 7'h47; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_647 = io_wen & io_addr[10:4] == 7'h47 ? io_wdata[20] : tag_regs_71[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_71 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_647; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_71 = _valid_to_be_T_644 ? io_wdata[19:0] : tag_regs_71[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_71_T = {valid_to_be_71,tag_to_be_71}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_653 = io_wen & io_addr[10:4] == 7'h48; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_656 = io_wen & io_addr[10:4] == 7'h48 ? io_wdata[20] : tag_regs_72[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_72 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_656; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_72 = _valid_to_be_T_653 ? io_wdata[19:0] : tag_regs_72[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_72_T = {valid_to_be_72,tag_to_be_72}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_662 = io_wen & io_addr[10:4] == 7'h49; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_665 = io_wen & io_addr[10:4] == 7'h49 ? io_wdata[20] : tag_regs_73[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_73 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_665; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_73 = _valid_to_be_T_662 ? io_wdata[19:0] : tag_regs_73[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_73_T = {valid_to_be_73,tag_to_be_73}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_671 = io_wen & io_addr[10:4] == 7'h4a; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_674 = io_wen & io_addr[10:4] == 7'h4a ? io_wdata[20] : tag_regs_74[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_74 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_674; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_74 = _valid_to_be_T_671 ? io_wdata[19:0] : tag_regs_74[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_74_T = {valid_to_be_74,tag_to_be_74}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_680 = io_wen & io_addr[10:4] == 7'h4b; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_683 = io_wen & io_addr[10:4] == 7'h4b ? io_wdata[20] : tag_regs_75[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_75 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_683; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_75 = _valid_to_be_T_680 ? io_wdata[19:0] : tag_regs_75[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_75_T = {valid_to_be_75,tag_to_be_75}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_689 = io_wen & io_addr[10:4] == 7'h4c; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_692 = io_wen & io_addr[10:4] == 7'h4c ? io_wdata[20] : tag_regs_76[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_76 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_692; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_76 = _valid_to_be_T_689 ? io_wdata[19:0] : tag_regs_76[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_76_T = {valid_to_be_76,tag_to_be_76}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_698 = io_wen & io_addr[10:4] == 7'h4d; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_701 = io_wen & io_addr[10:4] == 7'h4d ? io_wdata[20] : tag_regs_77[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_77 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_701; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_77 = _valid_to_be_T_698 ? io_wdata[19:0] : tag_regs_77[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_77_T = {valid_to_be_77,tag_to_be_77}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_707 = io_wen & io_addr[10:4] == 7'h4e; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_710 = io_wen & io_addr[10:4] == 7'h4e ? io_wdata[20] : tag_regs_78[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_78 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_710; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_78 = _valid_to_be_T_707 ? io_wdata[19:0] : tag_regs_78[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_78_T = {valid_to_be_78,tag_to_be_78}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_716 = io_wen & io_addr[10:4] == 7'h4f; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_719 = io_wen & io_addr[10:4] == 7'h4f ? io_wdata[20] : tag_regs_79[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_79 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_719; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_79 = _valid_to_be_T_716 ? io_wdata[19:0] : tag_regs_79[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_79_T = {valid_to_be_79,tag_to_be_79}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_725 = io_wen & io_addr[10:4] == 7'h50; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_728 = io_wen & io_addr[10:4] == 7'h50 ? io_wdata[20] : tag_regs_80[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_80 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_728; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_80 = _valid_to_be_T_725 ? io_wdata[19:0] : tag_regs_80[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_80_T = {valid_to_be_80,tag_to_be_80}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_734 = io_wen & io_addr[10:4] == 7'h51; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_737 = io_wen & io_addr[10:4] == 7'h51 ? io_wdata[20] : tag_regs_81[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_81 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_737; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_81 = _valid_to_be_T_734 ? io_wdata[19:0] : tag_regs_81[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_81_T = {valid_to_be_81,tag_to_be_81}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_743 = io_wen & io_addr[10:4] == 7'h52; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_746 = io_wen & io_addr[10:4] == 7'h52 ? io_wdata[20] : tag_regs_82[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_82 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_746; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_82 = _valid_to_be_T_743 ? io_wdata[19:0] : tag_regs_82[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_82_T = {valid_to_be_82,tag_to_be_82}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_752 = io_wen & io_addr[10:4] == 7'h53; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_755 = io_wen & io_addr[10:4] == 7'h53 ? io_wdata[20] : tag_regs_83[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_83 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_755; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_83 = _valid_to_be_T_752 ? io_wdata[19:0] : tag_regs_83[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_83_T = {valid_to_be_83,tag_to_be_83}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_761 = io_wen & io_addr[10:4] == 7'h54; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_764 = io_wen & io_addr[10:4] == 7'h54 ? io_wdata[20] : tag_regs_84[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_84 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_764; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_84 = _valid_to_be_T_761 ? io_wdata[19:0] : tag_regs_84[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_84_T = {valid_to_be_84,tag_to_be_84}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_770 = io_wen & io_addr[10:4] == 7'h55; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_773 = io_wen & io_addr[10:4] == 7'h55 ? io_wdata[20] : tag_regs_85[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_85 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_773; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_85 = _valid_to_be_T_770 ? io_wdata[19:0] : tag_regs_85[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_85_T = {valid_to_be_85,tag_to_be_85}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_779 = io_wen & io_addr[10:4] == 7'h56; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_782 = io_wen & io_addr[10:4] == 7'h56 ? io_wdata[20] : tag_regs_86[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_86 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_782; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_86 = _valid_to_be_T_779 ? io_wdata[19:0] : tag_regs_86[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_86_T = {valid_to_be_86,tag_to_be_86}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_788 = io_wen & io_addr[10:4] == 7'h57; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_791 = io_wen & io_addr[10:4] == 7'h57 ? io_wdata[20] : tag_regs_87[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_87 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_791; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_87 = _valid_to_be_T_788 ? io_wdata[19:0] : tag_regs_87[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_87_T = {valid_to_be_87,tag_to_be_87}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_797 = io_wen & io_addr[10:4] == 7'h58; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_800 = io_wen & io_addr[10:4] == 7'h58 ? io_wdata[20] : tag_regs_88[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_88 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_800; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_88 = _valid_to_be_T_797 ? io_wdata[19:0] : tag_regs_88[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_88_T = {valid_to_be_88,tag_to_be_88}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_806 = io_wen & io_addr[10:4] == 7'h59; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_809 = io_wen & io_addr[10:4] == 7'h59 ? io_wdata[20] : tag_regs_89[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_89 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_809; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_89 = _valid_to_be_T_806 ? io_wdata[19:0] : tag_regs_89[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_89_T = {valid_to_be_89,tag_to_be_89}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_815 = io_wen & io_addr[10:4] == 7'h5a; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_818 = io_wen & io_addr[10:4] == 7'h5a ? io_wdata[20] : tag_regs_90[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_90 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_818; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_90 = _valid_to_be_T_815 ? io_wdata[19:0] : tag_regs_90[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_90_T = {valid_to_be_90,tag_to_be_90}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_824 = io_wen & io_addr[10:4] == 7'h5b; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_827 = io_wen & io_addr[10:4] == 7'h5b ? io_wdata[20] : tag_regs_91[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_91 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_827; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_91 = _valid_to_be_T_824 ? io_wdata[19:0] : tag_regs_91[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_91_T = {valid_to_be_91,tag_to_be_91}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_833 = io_wen & io_addr[10:4] == 7'h5c; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_836 = io_wen & io_addr[10:4] == 7'h5c ? io_wdata[20] : tag_regs_92[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_92 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_836; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_92 = _valid_to_be_T_833 ? io_wdata[19:0] : tag_regs_92[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_92_T = {valid_to_be_92,tag_to_be_92}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_842 = io_wen & io_addr[10:4] == 7'h5d; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_845 = io_wen & io_addr[10:4] == 7'h5d ? io_wdata[20] : tag_regs_93[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_93 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_845; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_93 = _valid_to_be_T_842 ? io_wdata[19:0] : tag_regs_93[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_93_T = {valid_to_be_93,tag_to_be_93}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_851 = io_wen & io_addr[10:4] == 7'h5e; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_854 = io_wen & io_addr[10:4] == 7'h5e ? io_wdata[20] : tag_regs_94[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_94 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_854; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_94 = _valid_to_be_T_851 ? io_wdata[19:0] : tag_regs_94[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_94_T = {valid_to_be_94,tag_to_be_94}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_860 = io_wen & io_addr[10:4] == 7'h5f; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_863 = io_wen & io_addr[10:4] == 7'h5f ? io_wdata[20] : tag_regs_95[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_95 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_863; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_95 = _valid_to_be_T_860 ? io_wdata[19:0] : tag_regs_95[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_95_T = {valid_to_be_95,tag_to_be_95}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_869 = io_wen & io_addr[10:4] == 7'h60; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_872 = io_wen & io_addr[10:4] == 7'h60 ? io_wdata[20] : tag_regs_96[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_96 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_872; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_96 = _valid_to_be_T_869 ? io_wdata[19:0] : tag_regs_96[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_96_T = {valid_to_be_96,tag_to_be_96}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_878 = io_wen & io_addr[10:4] == 7'h61; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_881 = io_wen & io_addr[10:4] == 7'h61 ? io_wdata[20] : tag_regs_97[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_97 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_881; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_97 = _valid_to_be_T_878 ? io_wdata[19:0] : tag_regs_97[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_97_T = {valid_to_be_97,tag_to_be_97}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_887 = io_wen & io_addr[10:4] == 7'h62; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_890 = io_wen & io_addr[10:4] == 7'h62 ? io_wdata[20] : tag_regs_98[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_98 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_890; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_98 = _valid_to_be_T_887 ? io_wdata[19:0] : tag_regs_98[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_98_T = {valid_to_be_98,tag_to_be_98}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_896 = io_wen & io_addr[10:4] == 7'h63; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_899 = io_wen & io_addr[10:4] == 7'h63 ? io_wdata[20] : tag_regs_99[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_99 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_899; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_99 = _valid_to_be_T_896 ? io_wdata[19:0] : tag_regs_99[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_99_T = {valid_to_be_99,tag_to_be_99}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_905 = io_wen & io_addr[10:4] == 7'h64; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_908 = io_wen & io_addr[10:4] == 7'h64 ? io_wdata[20] : tag_regs_100[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_100 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_908; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_100 = _valid_to_be_T_905 ? io_wdata[19:0] : tag_regs_100[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_100_T = {valid_to_be_100,tag_to_be_100}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_914 = io_wen & io_addr[10:4] == 7'h65; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_917 = io_wen & io_addr[10:4] == 7'h65 ? io_wdata[20] : tag_regs_101[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_101 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_917; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_101 = _valid_to_be_T_914 ? io_wdata[19:0] : tag_regs_101[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_101_T = {valid_to_be_101,tag_to_be_101}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_923 = io_wen & io_addr[10:4] == 7'h66; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_926 = io_wen & io_addr[10:4] == 7'h66 ? io_wdata[20] : tag_regs_102[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_102 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_926; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_102 = _valid_to_be_T_923 ? io_wdata[19:0] : tag_regs_102[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_102_T = {valid_to_be_102,tag_to_be_102}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_932 = io_wen & io_addr[10:4] == 7'h67; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_935 = io_wen & io_addr[10:4] == 7'h67 ? io_wdata[20] : tag_regs_103[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_103 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_935; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_103 = _valid_to_be_T_932 ? io_wdata[19:0] : tag_regs_103[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_103_T = {valid_to_be_103,tag_to_be_103}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_941 = io_wen & io_addr[10:4] == 7'h68; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_944 = io_wen & io_addr[10:4] == 7'h68 ? io_wdata[20] : tag_regs_104[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_104 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_944; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_104 = _valid_to_be_T_941 ? io_wdata[19:0] : tag_regs_104[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_104_T = {valid_to_be_104,tag_to_be_104}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_950 = io_wen & io_addr[10:4] == 7'h69; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_953 = io_wen & io_addr[10:4] == 7'h69 ? io_wdata[20] : tag_regs_105[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_105 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_953; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_105 = _valid_to_be_T_950 ? io_wdata[19:0] : tag_regs_105[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_105_T = {valid_to_be_105,tag_to_be_105}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_959 = io_wen & io_addr[10:4] == 7'h6a; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_962 = io_wen & io_addr[10:4] == 7'h6a ? io_wdata[20] : tag_regs_106[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_106 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_962; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_106 = _valid_to_be_T_959 ? io_wdata[19:0] : tag_regs_106[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_106_T = {valid_to_be_106,tag_to_be_106}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_968 = io_wen & io_addr[10:4] == 7'h6b; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_971 = io_wen & io_addr[10:4] == 7'h6b ? io_wdata[20] : tag_regs_107[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_107 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_971; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_107 = _valid_to_be_T_968 ? io_wdata[19:0] : tag_regs_107[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_107_T = {valid_to_be_107,tag_to_be_107}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_977 = io_wen & io_addr[10:4] == 7'h6c; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_980 = io_wen & io_addr[10:4] == 7'h6c ? io_wdata[20] : tag_regs_108[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_108 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_980; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_108 = _valid_to_be_T_977 ? io_wdata[19:0] : tag_regs_108[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_108_T = {valid_to_be_108,tag_to_be_108}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_986 = io_wen & io_addr[10:4] == 7'h6d; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_989 = io_wen & io_addr[10:4] == 7'h6d ? io_wdata[20] : tag_regs_109[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_109 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_989; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_109 = _valid_to_be_T_986 ? io_wdata[19:0] : tag_regs_109[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_109_T = {valid_to_be_109,tag_to_be_109}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_995 = io_wen & io_addr[10:4] == 7'h6e; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_998 = io_wen & io_addr[10:4] == 7'h6e ? io_wdata[20] : tag_regs_110[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_110 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_998; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_110 = _valid_to_be_T_995 ? io_wdata[19:0] : tag_regs_110[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_110_T = {valid_to_be_110,tag_to_be_110}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1004 = io_wen & io_addr[10:4] == 7'h6f; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1007 = io_wen & io_addr[10:4] == 7'h6f ? io_wdata[20] : tag_regs_111[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_111 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1007; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_111 = _valid_to_be_T_1004 ? io_wdata[19:0] : tag_regs_111[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_111_T = {valid_to_be_111,tag_to_be_111}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1013 = io_wen & io_addr[10:4] == 7'h70; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1016 = io_wen & io_addr[10:4] == 7'h70 ? io_wdata[20] : tag_regs_112[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_112 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1016; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_112 = _valid_to_be_T_1013 ? io_wdata[19:0] : tag_regs_112[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_112_T = {valid_to_be_112,tag_to_be_112}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1022 = io_wen & io_addr[10:4] == 7'h71; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1025 = io_wen & io_addr[10:4] == 7'h71 ? io_wdata[20] : tag_regs_113[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_113 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1025; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_113 = _valid_to_be_T_1022 ? io_wdata[19:0] : tag_regs_113[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_113_T = {valid_to_be_113,tag_to_be_113}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1031 = io_wen & io_addr[10:4] == 7'h72; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1034 = io_wen & io_addr[10:4] == 7'h72 ? io_wdata[20] : tag_regs_114[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_114 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1034; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_114 = _valid_to_be_T_1031 ? io_wdata[19:0] : tag_regs_114[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_114_T = {valid_to_be_114,tag_to_be_114}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1040 = io_wen & io_addr[10:4] == 7'h73; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1043 = io_wen & io_addr[10:4] == 7'h73 ? io_wdata[20] : tag_regs_115[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_115 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1043; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_115 = _valid_to_be_T_1040 ? io_wdata[19:0] : tag_regs_115[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_115_T = {valid_to_be_115,tag_to_be_115}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1049 = io_wen & io_addr[10:4] == 7'h74; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1052 = io_wen & io_addr[10:4] == 7'h74 ? io_wdata[20] : tag_regs_116[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_116 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1052; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_116 = _valid_to_be_T_1049 ? io_wdata[19:0] : tag_regs_116[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_116_T = {valid_to_be_116,tag_to_be_116}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1058 = io_wen & io_addr[10:4] == 7'h75; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1061 = io_wen & io_addr[10:4] == 7'h75 ? io_wdata[20] : tag_regs_117[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_117 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1061; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_117 = _valid_to_be_T_1058 ? io_wdata[19:0] : tag_regs_117[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_117_T = {valid_to_be_117,tag_to_be_117}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1067 = io_wen & io_addr[10:4] == 7'h76; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1070 = io_wen & io_addr[10:4] == 7'h76 ? io_wdata[20] : tag_regs_118[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_118 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1070; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_118 = _valid_to_be_T_1067 ? io_wdata[19:0] : tag_regs_118[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_118_T = {valid_to_be_118,tag_to_be_118}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1076 = io_wen & io_addr[10:4] == 7'h77; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1079 = io_wen & io_addr[10:4] == 7'h77 ? io_wdata[20] : tag_regs_119[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_119 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1079; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_119 = _valid_to_be_T_1076 ? io_wdata[19:0] : tag_regs_119[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_119_T = {valid_to_be_119,tag_to_be_119}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1085 = io_wen & io_addr[10:4] == 7'h78; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1088 = io_wen & io_addr[10:4] == 7'h78 ? io_wdata[20] : tag_regs_120[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_120 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1088; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_120 = _valid_to_be_T_1085 ? io_wdata[19:0] : tag_regs_120[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_120_T = {valid_to_be_120,tag_to_be_120}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1094 = io_wen & io_addr[10:4] == 7'h79; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1097 = io_wen & io_addr[10:4] == 7'h79 ? io_wdata[20] : tag_regs_121[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_121 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1097; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_121 = _valid_to_be_T_1094 ? io_wdata[19:0] : tag_regs_121[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_121_T = {valid_to_be_121,tag_to_be_121}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1103 = io_wen & io_addr[10:4] == 7'h7a; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1106 = io_wen & io_addr[10:4] == 7'h7a ? io_wdata[20] : tag_regs_122[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_122 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1106; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_122 = _valid_to_be_T_1103 ? io_wdata[19:0] : tag_regs_122[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_122_T = {valid_to_be_122,tag_to_be_122}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1112 = io_wen & io_addr[10:4] == 7'h7b; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1115 = io_wen & io_addr[10:4] == 7'h7b ? io_wdata[20] : tag_regs_123[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_123 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1115; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_123 = _valid_to_be_T_1112 ? io_wdata[19:0] : tag_regs_123[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_123_T = {valid_to_be_123,tag_to_be_123}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1121 = io_wen & io_addr[10:4] == 7'h7c; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1124 = io_wen & io_addr[10:4] == 7'h7c ? io_wdata[20] : tag_regs_124[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_124 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1124; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_124 = _valid_to_be_T_1121 ? io_wdata[19:0] : tag_regs_124[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_124_T = {valid_to_be_124,tag_to_be_124}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1130 = io_wen & io_addr[10:4] == 7'h7d; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1133 = io_wen & io_addr[10:4] == 7'h7d ? io_wdata[20] : tag_regs_125[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_125 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1133; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_125 = _valid_to_be_T_1130 ? io_wdata[19:0] : tag_regs_125[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_125_T = {valid_to_be_125,tag_to_be_125}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1139 = io_wen & io_addr[10:4] == 7'h7e; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1142 = io_wen & io_addr[10:4] == 7'h7e ? io_wdata[20] : tag_regs_126[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_126 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1142; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_126 = _valid_to_be_T_1139 ? io_wdata[19:0] : tag_regs_126[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_126_T = {valid_to_be_126,tag_to_be_126}; // @[Cat.scala 31:58]
  wire  _valid_to_be_T_1148 = io_wen & io_addr[10:4] == 7'h7f; // @[icache_tag.scala 27:93]
  wire  _valid_to_be_T_1151 = io_wen & io_addr[10:4] == 7'h7f ? io_wdata[20] : tag_regs_127[20]; // @[icache_tag.scala 27:62]
  wire  valid_to_be_127 = io_tag_all_flush ? 1'h0 : _valid_to_be_T_1151; // @[icache_tag.scala 27:30]
  wire [19:0] tag_to_be_127 = _valid_to_be_T_1148 ? io_wdata[19:0] : tag_regs_127[19:0]; // @[icache_tag.scala 30:28]
  wire [20:0] _tag_regs_127_T = {valid_to_be_127,tag_to_be_127}; // @[Cat.scala 31:58]
  wire [7:0] _GEN_1 = 7'h1 == io_addr[10:4] ? tag_asid_regs_1 : tag_asid_regs_0; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_2 = 7'h2 == io_addr[10:4] ? tag_asid_regs_2 : _GEN_1; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_3 = 7'h3 == io_addr[10:4] ? tag_asid_regs_3 : _GEN_2; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_4 = 7'h4 == io_addr[10:4] ? tag_asid_regs_4 : _GEN_3; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_5 = 7'h5 == io_addr[10:4] ? tag_asid_regs_5 : _GEN_4; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_6 = 7'h6 == io_addr[10:4] ? tag_asid_regs_6 : _GEN_5; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_7 = 7'h7 == io_addr[10:4] ? tag_asid_regs_7 : _GEN_6; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_8 = 7'h8 == io_addr[10:4] ? tag_asid_regs_8 : _GEN_7; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_9 = 7'h9 == io_addr[10:4] ? tag_asid_regs_9 : _GEN_8; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_10 = 7'ha == io_addr[10:4] ? tag_asid_regs_10 : _GEN_9; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_11 = 7'hb == io_addr[10:4] ? tag_asid_regs_11 : _GEN_10; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_12 = 7'hc == io_addr[10:4] ? tag_asid_regs_12 : _GEN_11; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_13 = 7'hd == io_addr[10:4] ? tag_asid_regs_13 : _GEN_12; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_14 = 7'he == io_addr[10:4] ? tag_asid_regs_14 : _GEN_13; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_15 = 7'hf == io_addr[10:4] ? tag_asid_regs_15 : _GEN_14; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_16 = 7'h10 == io_addr[10:4] ? tag_asid_regs_16 : _GEN_15; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_17 = 7'h11 == io_addr[10:4] ? tag_asid_regs_17 : _GEN_16; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_18 = 7'h12 == io_addr[10:4] ? tag_asid_regs_18 : _GEN_17; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_19 = 7'h13 == io_addr[10:4] ? tag_asid_regs_19 : _GEN_18; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_20 = 7'h14 == io_addr[10:4] ? tag_asid_regs_20 : _GEN_19; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_21 = 7'h15 == io_addr[10:4] ? tag_asid_regs_21 : _GEN_20; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_22 = 7'h16 == io_addr[10:4] ? tag_asid_regs_22 : _GEN_21; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_23 = 7'h17 == io_addr[10:4] ? tag_asid_regs_23 : _GEN_22; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_24 = 7'h18 == io_addr[10:4] ? tag_asid_regs_24 : _GEN_23; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_25 = 7'h19 == io_addr[10:4] ? tag_asid_regs_25 : _GEN_24; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_26 = 7'h1a == io_addr[10:4] ? tag_asid_regs_26 : _GEN_25; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_27 = 7'h1b == io_addr[10:4] ? tag_asid_regs_27 : _GEN_26; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_28 = 7'h1c == io_addr[10:4] ? tag_asid_regs_28 : _GEN_27; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_29 = 7'h1d == io_addr[10:4] ? tag_asid_regs_29 : _GEN_28; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_30 = 7'h1e == io_addr[10:4] ? tag_asid_regs_30 : _GEN_29; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_31 = 7'h1f == io_addr[10:4] ? tag_asid_regs_31 : _GEN_30; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_32 = 7'h20 == io_addr[10:4] ? tag_asid_regs_32 : _GEN_31; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_33 = 7'h21 == io_addr[10:4] ? tag_asid_regs_33 : _GEN_32; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_34 = 7'h22 == io_addr[10:4] ? tag_asid_regs_34 : _GEN_33; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_35 = 7'h23 == io_addr[10:4] ? tag_asid_regs_35 : _GEN_34; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_36 = 7'h24 == io_addr[10:4] ? tag_asid_regs_36 : _GEN_35; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_37 = 7'h25 == io_addr[10:4] ? tag_asid_regs_37 : _GEN_36; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_38 = 7'h26 == io_addr[10:4] ? tag_asid_regs_38 : _GEN_37; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_39 = 7'h27 == io_addr[10:4] ? tag_asid_regs_39 : _GEN_38; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_40 = 7'h28 == io_addr[10:4] ? tag_asid_regs_40 : _GEN_39; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_41 = 7'h29 == io_addr[10:4] ? tag_asid_regs_41 : _GEN_40; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_42 = 7'h2a == io_addr[10:4] ? tag_asid_regs_42 : _GEN_41; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_43 = 7'h2b == io_addr[10:4] ? tag_asid_regs_43 : _GEN_42; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_44 = 7'h2c == io_addr[10:4] ? tag_asid_regs_44 : _GEN_43; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_45 = 7'h2d == io_addr[10:4] ? tag_asid_regs_45 : _GEN_44; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_46 = 7'h2e == io_addr[10:4] ? tag_asid_regs_46 : _GEN_45; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_47 = 7'h2f == io_addr[10:4] ? tag_asid_regs_47 : _GEN_46; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_48 = 7'h30 == io_addr[10:4] ? tag_asid_regs_48 : _GEN_47; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_49 = 7'h31 == io_addr[10:4] ? tag_asid_regs_49 : _GEN_48; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_50 = 7'h32 == io_addr[10:4] ? tag_asid_regs_50 : _GEN_49; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_51 = 7'h33 == io_addr[10:4] ? tag_asid_regs_51 : _GEN_50; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_52 = 7'h34 == io_addr[10:4] ? tag_asid_regs_52 : _GEN_51; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_53 = 7'h35 == io_addr[10:4] ? tag_asid_regs_53 : _GEN_52; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_54 = 7'h36 == io_addr[10:4] ? tag_asid_regs_54 : _GEN_53; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_55 = 7'h37 == io_addr[10:4] ? tag_asid_regs_55 : _GEN_54; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_56 = 7'h38 == io_addr[10:4] ? tag_asid_regs_56 : _GEN_55; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_57 = 7'h39 == io_addr[10:4] ? tag_asid_regs_57 : _GEN_56; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_58 = 7'h3a == io_addr[10:4] ? tag_asid_regs_58 : _GEN_57; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_59 = 7'h3b == io_addr[10:4] ? tag_asid_regs_59 : _GEN_58; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_60 = 7'h3c == io_addr[10:4] ? tag_asid_regs_60 : _GEN_59; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_61 = 7'h3d == io_addr[10:4] ? tag_asid_regs_61 : _GEN_60; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_62 = 7'h3e == io_addr[10:4] ? tag_asid_regs_62 : _GEN_61; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_63 = 7'h3f == io_addr[10:4] ? tag_asid_regs_63 : _GEN_62; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_64 = 7'h40 == io_addr[10:4] ? tag_asid_regs_64 : _GEN_63; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_65 = 7'h41 == io_addr[10:4] ? tag_asid_regs_65 : _GEN_64; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_66 = 7'h42 == io_addr[10:4] ? tag_asid_regs_66 : _GEN_65; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_67 = 7'h43 == io_addr[10:4] ? tag_asid_regs_67 : _GEN_66; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_68 = 7'h44 == io_addr[10:4] ? tag_asid_regs_68 : _GEN_67; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_69 = 7'h45 == io_addr[10:4] ? tag_asid_regs_69 : _GEN_68; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_70 = 7'h46 == io_addr[10:4] ? tag_asid_regs_70 : _GEN_69; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_71 = 7'h47 == io_addr[10:4] ? tag_asid_regs_71 : _GEN_70; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_72 = 7'h48 == io_addr[10:4] ? tag_asid_regs_72 : _GEN_71; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_73 = 7'h49 == io_addr[10:4] ? tag_asid_regs_73 : _GEN_72; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_74 = 7'h4a == io_addr[10:4] ? tag_asid_regs_74 : _GEN_73; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_75 = 7'h4b == io_addr[10:4] ? tag_asid_regs_75 : _GEN_74; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_76 = 7'h4c == io_addr[10:4] ? tag_asid_regs_76 : _GEN_75; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_77 = 7'h4d == io_addr[10:4] ? tag_asid_regs_77 : _GEN_76; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_78 = 7'h4e == io_addr[10:4] ? tag_asid_regs_78 : _GEN_77; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_79 = 7'h4f == io_addr[10:4] ? tag_asid_regs_79 : _GEN_78; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_80 = 7'h50 == io_addr[10:4] ? tag_asid_regs_80 : _GEN_79; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_81 = 7'h51 == io_addr[10:4] ? tag_asid_regs_81 : _GEN_80; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_82 = 7'h52 == io_addr[10:4] ? tag_asid_regs_82 : _GEN_81; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_83 = 7'h53 == io_addr[10:4] ? tag_asid_regs_83 : _GEN_82; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_84 = 7'h54 == io_addr[10:4] ? tag_asid_regs_84 : _GEN_83; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_85 = 7'h55 == io_addr[10:4] ? tag_asid_regs_85 : _GEN_84; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_86 = 7'h56 == io_addr[10:4] ? tag_asid_regs_86 : _GEN_85; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_87 = 7'h57 == io_addr[10:4] ? tag_asid_regs_87 : _GEN_86; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_88 = 7'h58 == io_addr[10:4] ? tag_asid_regs_88 : _GEN_87; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_89 = 7'h59 == io_addr[10:4] ? tag_asid_regs_89 : _GEN_88; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_90 = 7'h5a == io_addr[10:4] ? tag_asid_regs_90 : _GEN_89; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_91 = 7'h5b == io_addr[10:4] ? tag_asid_regs_91 : _GEN_90; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_92 = 7'h5c == io_addr[10:4] ? tag_asid_regs_92 : _GEN_91; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_93 = 7'h5d == io_addr[10:4] ? tag_asid_regs_93 : _GEN_92; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_94 = 7'h5e == io_addr[10:4] ? tag_asid_regs_94 : _GEN_93; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_95 = 7'h5f == io_addr[10:4] ? tag_asid_regs_95 : _GEN_94; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_96 = 7'h60 == io_addr[10:4] ? tag_asid_regs_96 : _GEN_95; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_97 = 7'h61 == io_addr[10:4] ? tag_asid_regs_97 : _GEN_96; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_98 = 7'h62 == io_addr[10:4] ? tag_asid_regs_98 : _GEN_97; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_99 = 7'h63 == io_addr[10:4] ? tag_asid_regs_99 : _GEN_98; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_100 = 7'h64 == io_addr[10:4] ? tag_asid_regs_100 : _GEN_99; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_101 = 7'h65 == io_addr[10:4] ? tag_asid_regs_101 : _GEN_100; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_102 = 7'h66 == io_addr[10:4] ? tag_asid_regs_102 : _GEN_101; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_103 = 7'h67 == io_addr[10:4] ? tag_asid_regs_103 : _GEN_102; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_104 = 7'h68 == io_addr[10:4] ? tag_asid_regs_104 : _GEN_103; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_105 = 7'h69 == io_addr[10:4] ? tag_asid_regs_105 : _GEN_104; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_106 = 7'h6a == io_addr[10:4] ? tag_asid_regs_106 : _GEN_105; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_107 = 7'h6b == io_addr[10:4] ? tag_asid_regs_107 : _GEN_106; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_108 = 7'h6c == io_addr[10:4] ? tag_asid_regs_108 : _GEN_107; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_109 = 7'h6d == io_addr[10:4] ? tag_asid_regs_109 : _GEN_108; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_110 = 7'h6e == io_addr[10:4] ? tag_asid_regs_110 : _GEN_109; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_111 = 7'h6f == io_addr[10:4] ? tag_asid_regs_111 : _GEN_110; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_112 = 7'h70 == io_addr[10:4] ? tag_asid_regs_112 : _GEN_111; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_113 = 7'h71 == io_addr[10:4] ? tag_asid_regs_113 : _GEN_112; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_114 = 7'h72 == io_addr[10:4] ? tag_asid_regs_114 : _GEN_113; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_115 = 7'h73 == io_addr[10:4] ? tag_asid_regs_115 : _GEN_114; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_116 = 7'h74 == io_addr[10:4] ? tag_asid_regs_116 : _GEN_115; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_117 = 7'h75 == io_addr[10:4] ? tag_asid_regs_117 : _GEN_116; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_118 = 7'h76 == io_addr[10:4] ? tag_asid_regs_118 : _GEN_117; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_119 = 7'h77 == io_addr[10:4] ? tag_asid_regs_119 : _GEN_118; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_120 = 7'h78 == io_addr[10:4] ? tag_asid_regs_120 : _GEN_119; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_121 = 7'h79 == io_addr[10:4] ? tag_asid_regs_121 : _GEN_120; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_122 = 7'h7a == io_addr[10:4] ? tag_asid_regs_122 : _GEN_121; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_123 = 7'h7b == io_addr[10:4] ? tag_asid_regs_123 : _GEN_122; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_124 = 7'h7c == io_addr[10:4] ? tag_asid_regs_124 : _GEN_123; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_125 = 7'h7d == io_addr[10:4] ? tag_asid_regs_125 : _GEN_124; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_126 = 7'h7e == io_addr[10:4] ? tag_asid_regs_126 : _GEN_125; // @[icache_tag.scala 33:{40,40}]
  wire [7:0] _GEN_127 = 7'h7f == io_addr[10:4] ? tag_asid_regs_127 : _GEN_126; // @[icache_tag.scala 33:{40,40}]
  wire [21:0] _GEN_257 = 7'h1 == io_addr[10:4] ? tag_regs_1 : tag_regs_0; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_258 = 7'h2 == io_addr[10:4] ? tag_regs_2 : _GEN_257; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_259 = 7'h3 == io_addr[10:4] ? tag_regs_3 : _GEN_258; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_260 = 7'h4 == io_addr[10:4] ? tag_regs_4 : _GEN_259; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_261 = 7'h5 == io_addr[10:4] ? tag_regs_5 : _GEN_260; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_262 = 7'h6 == io_addr[10:4] ? tag_regs_6 : _GEN_261; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_263 = 7'h7 == io_addr[10:4] ? tag_regs_7 : _GEN_262; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_264 = 7'h8 == io_addr[10:4] ? tag_regs_8 : _GEN_263; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_265 = 7'h9 == io_addr[10:4] ? tag_regs_9 : _GEN_264; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_266 = 7'ha == io_addr[10:4] ? tag_regs_10 : _GEN_265; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_267 = 7'hb == io_addr[10:4] ? tag_regs_11 : _GEN_266; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_268 = 7'hc == io_addr[10:4] ? tag_regs_12 : _GEN_267; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_269 = 7'hd == io_addr[10:4] ? tag_regs_13 : _GEN_268; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_270 = 7'he == io_addr[10:4] ? tag_regs_14 : _GEN_269; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_271 = 7'hf == io_addr[10:4] ? tag_regs_15 : _GEN_270; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_272 = 7'h10 == io_addr[10:4] ? tag_regs_16 : _GEN_271; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_273 = 7'h11 == io_addr[10:4] ? tag_regs_17 : _GEN_272; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_274 = 7'h12 == io_addr[10:4] ? tag_regs_18 : _GEN_273; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_275 = 7'h13 == io_addr[10:4] ? tag_regs_19 : _GEN_274; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_276 = 7'h14 == io_addr[10:4] ? tag_regs_20 : _GEN_275; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_277 = 7'h15 == io_addr[10:4] ? tag_regs_21 : _GEN_276; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_278 = 7'h16 == io_addr[10:4] ? tag_regs_22 : _GEN_277; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_279 = 7'h17 == io_addr[10:4] ? tag_regs_23 : _GEN_278; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_280 = 7'h18 == io_addr[10:4] ? tag_regs_24 : _GEN_279; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_281 = 7'h19 == io_addr[10:4] ? tag_regs_25 : _GEN_280; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_282 = 7'h1a == io_addr[10:4] ? tag_regs_26 : _GEN_281; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_283 = 7'h1b == io_addr[10:4] ? tag_regs_27 : _GEN_282; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_284 = 7'h1c == io_addr[10:4] ? tag_regs_28 : _GEN_283; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_285 = 7'h1d == io_addr[10:4] ? tag_regs_29 : _GEN_284; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_286 = 7'h1e == io_addr[10:4] ? tag_regs_30 : _GEN_285; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_287 = 7'h1f == io_addr[10:4] ? tag_regs_31 : _GEN_286; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_288 = 7'h20 == io_addr[10:4] ? tag_regs_32 : _GEN_287; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_289 = 7'h21 == io_addr[10:4] ? tag_regs_33 : _GEN_288; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_290 = 7'h22 == io_addr[10:4] ? tag_regs_34 : _GEN_289; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_291 = 7'h23 == io_addr[10:4] ? tag_regs_35 : _GEN_290; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_292 = 7'h24 == io_addr[10:4] ? tag_regs_36 : _GEN_291; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_293 = 7'h25 == io_addr[10:4] ? tag_regs_37 : _GEN_292; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_294 = 7'h26 == io_addr[10:4] ? tag_regs_38 : _GEN_293; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_295 = 7'h27 == io_addr[10:4] ? tag_regs_39 : _GEN_294; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_296 = 7'h28 == io_addr[10:4] ? tag_regs_40 : _GEN_295; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_297 = 7'h29 == io_addr[10:4] ? tag_regs_41 : _GEN_296; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_298 = 7'h2a == io_addr[10:4] ? tag_regs_42 : _GEN_297; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_299 = 7'h2b == io_addr[10:4] ? tag_regs_43 : _GEN_298; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_300 = 7'h2c == io_addr[10:4] ? tag_regs_44 : _GEN_299; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_301 = 7'h2d == io_addr[10:4] ? tag_regs_45 : _GEN_300; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_302 = 7'h2e == io_addr[10:4] ? tag_regs_46 : _GEN_301; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_303 = 7'h2f == io_addr[10:4] ? tag_regs_47 : _GEN_302; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_304 = 7'h30 == io_addr[10:4] ? tag_regs_48 : _GEN_303; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_305 = 7'h31 == io_addr[10:4] ? tag_regs_49 : _GEN_304; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_306 = 7'h32 == io_addr[10:4] ? tag_regs_50 : _GEN_305; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_307 = 7'h33 == io_addr[10:4] ? tag_regs_51 : _GEN_306; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_308 = 7'h34 == io_addr[10:4] ? tag_regs_52 : _GEN_307; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_309 = 7'h35 == io_addr[10:4] ? tag_regs_53 : _GEN_308; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_310 = 7'h36 == io_addr[10:4] ? tag_regs_54 : _GEN_309; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_311 = 7'h37 == io_addr[10:4] ? tag_regs_55 : _GEN_310; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_312 = 7'h38 == io_addr[10:4] ? tag_regs_56 : _GEN_311; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_313 = 7'h39 == io_addr[10:4] ? tag_regs_57 : _GEN_312; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_314 = 7'h3a == io_addr[10:4] ? tag_regs_58 : _GEN_313; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_315 = 7'h3b == io_addr[10:4] ? tag_regs_59 : _GEN_314; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_316 = 7'h3c == io_addr[10:4] ? tag_regs_60 : _GEN_315; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_317 = 7'h3d == io_addr[10:4] ? tag_regs_61 : _GEN_316; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_318 = 7'h3e == io_addr[10:4] ? tag_regs_62 : _GEN_317; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_319 = 7'h3f == io_addr[10:4] ? tag_regs_63 : _GEN_318; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_320 = 7'h40 == io_addr[10:4] ? tag_regs_64 : _GEN_319; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_321 = 7'h41 == io_addr[10:4] ? tag_regs_65 : _GEN_320; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_322 = 7'h42 == io_addr[10:4] ? tag_regs_66 : _GEN_321; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_323 = 7'h43 == io_addr[10:4] ? tag_regs_67 : _GEN_322; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_324 = 7'h44 == io_addr[10:4] ? tag_regs_68 : _GEN_323; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_325 = 7'h45 == io_addr[10:4] ? tag_regs_69 : _GEN_324; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_326 = 7'h46 == io_addr[10:4] ? tag_regs_70 : _GEN_325; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_327 = 7'h47 == io_addr[10:4] ? tag_regs_71 : _GEN_326; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_328 = 7'h48 == io_addr[10:4] ? tag_regs_72 : _GEN_327; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_329 = 7'h49 == io_addr[10:4] ? tag_regs_73 : _GEN_328; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_330 = 7'h4a == io_addr[10:4] ? tag_regs_74 : _GEN_329; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_331 = 7'h4b == io_addr[10:4] ? tag_regs_75 : _GEN_330; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_332 = 7'h4c == io_addr[10:4] ? tag_regs_76 : _GEN_331; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_333 = 7'h4d == io_addr[10:4] ? tag_regs_77 : _GEN_332; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_334 = 7'h4e == io_addr[10:4] ? tag_regs_78 : _GEN_333; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_335 = 7'h4f == io_addr[10:4] ? tag_regs_79 : _GEN_334; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_336 = 7'h50 == io_addr[10:4] ? tag_regs_80 : _GEN_335; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_337 = 7'h51 == io_addr[10:4] ? tag_regs_81 : _GEN_336; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_338 = 7'h52 == io_addr[10:4] ? tag_regs_82 : _GEN_337; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_339 = 7'h53 == io_addr[10:4] ? tag_regs_83 : _GEN_338; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_340 = 7'h54 == io_addr[10:4] ? tag_regs_84 : _GEN_339; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_341 = 7'h55 == io_addr[10:4] ? tag_regs_85 : _GEN_340; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_342 = 7'h56 == io_addr[10:4] ? tag_regs_86 : _GEN_341; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_343 = 7'h57 == io_addr[10:4] ? tag_regs_87 : _GEN_342; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_344 = 7'h58 == io_addr[10:4] ? tag_regs_88 : _GEN_343; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_345 = 7'h59 == io_addr[10:4] ? tag_regs_89 : _GEN_344; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_346 = 7'h5a == io_addr[10:4] ? tag_regs_90 : _GEN_345; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_347 = 7'h5b == io_addr[10:4] ? tag_regs_91 : _GEN_346; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_348 = 7'h5c == io_addr[10:4] ? tag_regs_92 : _GEN_347; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_349 = 7'h5d == io_addr[10:4] ? tag_regs_93 : _GEN_348; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_350 = 7'h5e == io_addr[10:4] ? tag_regs_94 : _GEN_349; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_351 = 7'h5f == io_addr[10:4] ? tag_regs_95 : _GEN_350; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_352 = 7'h60 == io_addr[10:4] ? tag_regs_96 : _GEN_351; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_353 = 7'h61 == io_addr[10:4] ? tag_regs_97 : _GEN_352; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_354 = 7'h62 == io_addr[10:4] ? tag_regs_98 : _GEN_353; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_355 = 7'h63 == io_addr[10:4] ? tag_regs_99 : _GEN_354; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_356 = 7'h64 == io_addr[10:4] ? tag_regs_100 : _GEN_355; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_357 = 7'h65 == io_addr[10:4] ? tag_regs_101 : _GEN_356; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_358 = 7'h66 == io_addr[10:4] ? tag_regs_102 : _GEN_357; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_359 = 7'h67 == io_addr[10:4] ? tag_regs_103 : _GEN_358; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_360 = 7'h68 == io_addr[10:4] ? tag_regs_104 : _GEN_359; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_361 = 7'h69 == io_addr[10:4] ? tag_regs_105 : _GEN_360; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_362 = 7'h6a == io_addr[10:4] ? tag_regs_106 : _GEN_361; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_363 = 7'h6b == io_addr[10:4] ? tag_regs_107 : _GEN_362; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_364 = 7'h6c == io_addr[10:4] ? tag_regs_108 : _GEN_363; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_365 = 7'h6d == io_addr[10:4] ? tag_regs_109 : _GEN_364; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_366 = 7'h6e == io_addr[10:4] ? tag_regs_110 : _GEN_365; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_367 = 7'h6f == io_addr[10:4] ? tag_regs_111 : _GEN_366; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_368 = 7'h70 == io_addr[10:4] ? tag_regs_112 : _GEN_367; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_369 = 7'h71 == io_addr[10:4] ? tag_regs_113 : _GEN_368; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_370 = 7'h72 == io_addr[10:4] ? tag_regs_114 : _GEN_369; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_371 = 7'h73 == io_addr[10:4] ? tag_regs_115 : _GEN_370; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_372 = 7'h74 == io_addr[10:4] ? tag_regs_116 : _GEN_371; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_373 = 7'h75 == io_addr[10:4] ? tag_regs_117 : _GEN_372; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_374 = 7'h76 == io_addr[10:4] ? tag_regs_118 : _GEN_373; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_375 = 7'h77 == io_addr[10:4] ? tag_regs_119 : _GEN_374; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_376 = 7'h78 == io_addr[10:4] ? tag_regs_120 : _GEN_375; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_377 = 7'h79 == io_addr[10:4] ? tag_regs_121 : _GEN_376; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_378 = 7'h7a == io_addr[10:4] ? tag_regs_122 : _GEN_377; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_379 = 7'h7b == io_addr[10:4] ? tag_regs_123 : _GEN_378; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_380 = 7'h7c == io_addr[10:4] ? tag_regs_124 : _GEN_379; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_381 = 7'h7d == io_addr[10:4] ? tag_regs_125 : _GEN_380; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_382 = 7'h7e == io_addr[10:4] ? tag_regs_126 : _GEN_381; // @[icache_tag.scala 36:{22,22}]
  wire [21:0] _GEN_383 = 7'h7f == io_addr[10:4] ? tag_regs_127 : _GEN_382; // @[icache_tag.scala 36:{22,22}]
  assign io_hit = _GEN_383[20:0] == io_addr[31:11] & _GEN_127 == 8'h0; // @[icache_tag.scala 37:50]
  assign io_valid = _GEN_383[20]; // @[icache_tag.scala 36:22]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_0 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_0 <= {{1'd0}, _tag_regs_0_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_1 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_1 <= {{1'd0}, _tag_regs_1_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_2 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_2 <= {{1'd0}, _tag_regs_2_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_3 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_3 <= {{1'd0}, _tag_regs_3_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_4 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_4 <= {{1'd0}, _tag_regs_4_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_5 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_5 <= {{1'd0}, _tag_regs_5_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_6 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_6 <= {{1'd0}, _tag_regs_6_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_7 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_7 <= {{1'd0}, _tag_regs_7_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_8 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_8 <= {{1'd0}, _tag_regs_8_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_9 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_9 <= {{1'd0}, _tag_regs_9_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_10 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_10 <= {{1'd0}, _tag_regs_10_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_11 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_11 <= {{1'd0}, _tag_regs_11_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_12 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_12 <= {{1'd0}, _tag_regs_12_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_13 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_13 <= {{1'd0}, _tag_regs_13_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_14 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_14 <= {{1'd0}, _tag_regs_14_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_15 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_15 <= {{1'd0}, _tag_regs_15_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_16 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_16 <= {{1'd0}, _tag_regs_16_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_17 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_17 <= {{1'd0}, _tag_regs_17_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_18 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_18 <= {{1'd0}, _tag_regs_18_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_19 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_19 <= {{1'd0}, _tag_regs_19_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_20 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_20 <= {{1'd0}, _tag_regs_20_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_21 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_21 <= {{1'd0}, _tag_regs_21_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_22 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_22 <= {{1'd0}, _tag_regs_22_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_23 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_23 <= {{1'd0}, _tag_regs_23_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_24 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_24 <= {{1'd0}, _tag_regs_24_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_25 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_25 <= {{1'd0}, _tag_regs_25_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_26 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_26 <= {{1'd0}, _tag_regs_26_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_27 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_27 <= {{1'd0}, _tag_regs_27_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_28 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_28 <= {{1'd0}, _tag_regs_28_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_29 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_29 <= {{1'd0}, _tag_regs_29_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_30 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_30 <= {{1'd0}, _tag_regs_30_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_31 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_31 <= {{1'd0}, _tag_regs_31_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_32 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_32 <= {{1'd0}, _tag_regs_32_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_33 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_33 <= {{1'd0}, _tag_regs_33_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_34 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_34 <= {{1'd0}, _tag_regs_34_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_35 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_35 <= {{1'd0}, _tag_regs_35_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_36 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_36 <= {{1'd0}, _tag_regs_36_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_37 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_37 <= {{1'd0}, _tag_regs_37_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_38 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_38 <= {{1'd0}, _tag_regs_38_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_39 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_39 <= {{1'd0}, _tag_regs_39_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_40 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_40 <= {{1'd0}, _tag_regs_40_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_41 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_41 <= {{1'd0}, _tag_regs_41_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_42 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_42 <= {{1'd0}, _tag_regs_42_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_43 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_43 <= {{1'd0}, _tag_regs_43_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_44 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_44 <= {{1'd0}, _tag_regs_44_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_45 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_45 <= {{1'd0}, _tag_regs_45_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_46 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_46 <= {{1'd0}, _tag_regs_46_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_47 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_47 <= {{1'd0}, _tag_regs_47_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_48 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_48 <= {{1'd0}, _tag_regs_48_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_49 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_49 <= {{1'd0}, _tag_regs_49_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_50 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_50 <= {{1'd0}, _tag_regs_50_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_51 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_51 <= {{1'd0}, _tag_regs_51_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_52 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_52 <= {{1'd0}, _tag_regs_52_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_53 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_53 <= {{1'd0}, _tag_regs_53_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_54 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_54 <= {{1'd0}, _tag_regs_54_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_55 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_55 <= {{1'd0}, _tag_regs_55_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_56 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_56 <= {{1'd0}, _tag_regs_56_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_57 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_57 <= {{1'd0}, _tag_regs_57_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_58 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_58 <= {{1'd0}, _tag_regs_58_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_59 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_59 <= {{1'd0}, _tag_regs_59_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_60 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_60 <= {{1'd0}, _tag_regs_60_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_61 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_61 <= {{1'd0}, _tag_regs_61_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_62 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_62 <= {{1'd0}, _tag_regs_62_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_63 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_63 <= {{1'd0}, _tag_regs_63_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_64 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_64 <= {{1'd0}, _tag_regs_64_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_65 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_65 <= {{1'd0}, _tag_regs_65_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_66 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_66 <= {{1'd0}, _tag_regs_66_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_67 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_67 <= {{1'd0}, _tag_regs_67_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_68 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_68 <= {{1'd0}, _tag_regs_68_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_69 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_69 <= {{1'd0}, _tag_regs_69_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_70 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_70 <= {{1'd0}, _tag_regs_70_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_71 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_71 <= {{1'd0}, _tag_regs_71_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_72 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_72 <= {{1'd0}, _tag_regs_72_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_73 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_73 <= {{1'd0}, _tag_regs_73_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_74 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_74 <= {{1'd0}, _tag_regs_74_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_75 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_75 <= {{1'd0}, _tag_regs_75_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_76 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_76 <= {{1'd0}, _tag_regs_76_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_77 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_77 <= {{1'd0}, _tag_regs_77_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_78 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_78 <= {{1'd0}, _tag_regs_78_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_79 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_79 <= {{1'd0}, _tag_regs_79_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_80 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_80 <= {{1'd0}, _tag_regs_80_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_81 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_81 <= {{1'd0}, _tag_regs_81_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_82 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_82 <= {{1'd0}, _tag_regs_82_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_83 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_83 <= {{1'd0}, _tag_regs_83_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_84 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_84 <= {{1'd0}, _tag_regs_84_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_85 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_85 <= {{1'd0}, _tag_regs_85_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_86 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_86 <= {{1'd0}, _tag_regs_86_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_87 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_87 <= {{1'd0}, _tag_regs_87_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_88 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_88 <= {{1'd0}, _tag_regs_88_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_89 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_89 <= {{1'd0}, _tag_regs_89_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_90 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_90 <= {{1'd0}, _tag_regs_90_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_91 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_91 <= {{1'd0}, _tag_regs_91_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_92 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_92 <= {{1'd0}, _tag_regs_92_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_93 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_93 <= {{1'd0}, _tag_regs_93_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_94 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_94 <= {{1'd0}, _tag_regs_94_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_95 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_95 <= {{1'd0}, _tag_regs_95_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_96 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_96 <= {{1'd0}, _tag_regs_96_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_97 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_97 <= {{1'd0}, _tag_regs_97_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_98 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_98 <= {{1'd0}, _tag_regs_98_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_99 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_99 <= {{1'd0}, _tag_regs_99_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_100 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_100 <= {{1'd0}, _tag_regs_100_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_101 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_101 <= {{1'd0}, _tag_regs_101_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_102 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_102 <= {{1'd0}, _tag_regs_102_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_103 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_103 <= {{1'd0}, _tag_regs_103_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_104 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_104 <= {{1'd0}, _tag_regs_104_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_105 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_105 <= {{1'd0}, _tag_regs_105_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_106 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_106 <= {{1'd0}, _tag_regs_106_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_107 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_107 <= {{1'd0}, _tag_regs_107_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_108 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_108 <= {{1'd0}, _tag_regs_108_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_109 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_109 <= {{1'd0}, _tag_regs_109_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_110 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_110 <= {{1'd0}, _tag_regs_110_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_111 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_111 <= {{1'd0}, _tag_regs_111_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_112 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_112 <= {{1'd0}, _tag_regs_112_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_113 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_113 <= {{1'd0}, _tag_regs_113_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_114 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_114 <= {{1'd0}, _tag_regs_114_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_115 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_115 <= {{1'd0}, _tag_regs_115_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_116 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_116 <= {{1'd0}, _tag_regs_116_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_117 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_117 <= {{1'd0}, _tag_regs_117_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_118 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_118 <= {{1'd0}, _tag_regs_118_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_119 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_119 <= {{1'd0}, _tag_regs_119_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_120 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_120 <= {{1'd0}, _tag_regs_120_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_121 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_121 <= {{1'd0}, _tag_regs_121_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_122 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_122 <= {{1'd0}, _tag_regs_122_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_123 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_123 <= {{1'd0}, _tag_regs_123_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_124 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_124 <= {{1'd0}, _tag_regs_124_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_125 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_125 <= {{1'd0}, _tag_regs_125_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_126 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_126 <= {{1'd0}, _tag_regs_126_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 21:27]
      tag_regs_127 <= 22'h0; // @[icache_tag.scala 21:27]
    end else begin
      tag_regs_127 <= {{1'd0}, _tag_regs_127_T}; // @[icache_tag.scala 31:25]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_0 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h0 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_0 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_0 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_0 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_0 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_1 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h1 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_1 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_1 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_1 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_1 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_2 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h2 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_2 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_2 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_2 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_2 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_3 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h3 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_3 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_3 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_3 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_3 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_4 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h4 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_4 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_4 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_4 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_4 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_5 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h5 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_5 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_5 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_5 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_5 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_6 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h6 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_6 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_6 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_6 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_6 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_7 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h7 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_7 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_7 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_7 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_7 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_8 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h8 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_8 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_8 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_8 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_8 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_9 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h9 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_9 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_9 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_9 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_9 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_10 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'ha == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_10 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_10 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_10 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_10 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_11 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'hb == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_11 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_11 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_11 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_11 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_12 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'hc == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_12 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_12 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_12 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_12 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_13 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'hd == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_13 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_13 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_13 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_13 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_14 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'he == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_14 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_14 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_14 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_14 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_15 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'hf == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_15 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_15 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_15 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_15 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_16 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h10 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_16 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_16 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_16 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_16 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_17 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h11 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_17 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_17 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_17 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_17 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_18 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h12 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_18 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_18 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_18 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_18 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_19 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h13 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_19 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_19 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_19 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_19 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_20 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h14 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_20 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_20 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_20 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_20 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_21 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h15 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_21 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_21 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_21 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_21 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_22 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h16 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_22 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_22 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_22 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_22 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_23 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h17 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_23 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_23 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_23 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_23 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_24 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h18 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_24 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_24 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_24 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_24 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_25 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h19 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_25 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_25 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_25 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_25 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_26 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h1a == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_26 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_26 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_26 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_26 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_27 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h1b == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_27 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_27 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_27 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_27 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_28 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h1c == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_28 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_28 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_28 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_28 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_29 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h1d == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_29 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_29 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_29 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_29 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_30 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h1e == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_30 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_30 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_30 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_30 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_31 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h1f == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_31 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_31 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_31 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_31 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_32 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h20 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_32 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_32 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_32 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_32 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_33 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h21 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_33 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_33 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_33 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_33 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_34 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h22 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_34 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_34 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_34 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_34 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_35 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h23 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_35 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_35 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_35 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_35 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_36 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h24 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_36 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_36 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_36 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_36 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_37 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h25 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_37 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_37 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_37 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_37 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_38 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h26 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_38 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_38 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_38 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_38 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_39 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h27 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_39 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_39 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_39 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_39 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_40 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h28 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_40 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_40 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_40 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_40 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_41 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h29 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_41 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_41 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_41 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_41 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_42 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h2a == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_42 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_42 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_42 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_42 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_43 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h2b == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_43 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_43 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_43 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_43 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_44 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h2c == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_44 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_44 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_44 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_44 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_45 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h2d == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_45 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_45 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_45 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_45 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_46 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h2e == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_46 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_46 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_46 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_46 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_47 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h2f == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_47 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_47 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_47 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_47 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_48 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h30 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_48 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_48 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_48 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_48 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_49 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h31 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_49 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_49 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_49 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_49 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_50 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h32 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_50 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_50 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_50 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_50 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_51 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h33 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_51 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_51 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_51 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_51 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_52 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h34 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_52 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_52 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_52 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_52 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_53 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h35 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_53 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_53 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_53 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_53 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_54 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h36 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_54 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_54 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_54 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_54 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_55 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h37 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_55 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_55 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_55 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_55 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_56 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h38 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_56 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_56 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_56 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_56 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_57 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h39 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_57 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_57 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_57 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_57 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_58 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h3a == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_58 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_58 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_58 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_58 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_59 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h3b == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_59 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_59 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_59 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_59 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_60 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h3c == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_60 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_60 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_60 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_60 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_61 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h3d == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_61 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_61 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_61 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_61 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_62 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h3e == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_62 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_62 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_62 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_62 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_63 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h3f == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_63 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_63 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_63 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_63 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_64 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h40 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_64 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_64 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_64 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_64 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_65 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h41 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_65 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_65 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_65 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_65 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_66 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h42 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_66 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_66 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_66 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_66 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_67 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h43 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_67 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_67 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_67 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_67 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_68 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h44 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_68 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_68 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_68 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_68 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_69 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h45 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_69 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_69 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_69 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_69 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_70 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h46 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_70 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_70 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_70 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_70 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_71 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h47 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_71 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_71 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_71 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_71 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_72 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h48 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_72 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_72 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_72 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_72 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_73 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h49 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_73 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_73 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_73 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_73 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_74 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h4a == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_74 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_74 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_74 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_74 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_75 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h4b == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_75 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_75 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_75 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_75 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_76 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h4c == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_76 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_76 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_76 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_76 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_77 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h4d == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_77 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_77 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_77 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_77 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_78 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h4e == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_78 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_78 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_78 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_78 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_79 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h4f == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_79 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_79 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_79 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_79 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_80 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h50 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_80 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_80 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_80 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_80 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_81 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h51 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_81 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_81 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_81 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_81 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_82 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h52 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_82 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_82 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_82 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_82 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_83 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h53 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_83 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_83 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_83 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_83 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_84 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h54 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_84 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_84 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_84 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_84 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_85 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h55 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_85 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_85 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_85 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_85 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_86 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h56 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_86 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_86 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_86 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_86 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_87 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h57 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_87 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_87 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_87 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_87 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_88 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h58 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_88 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_88 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_88 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_88 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_89 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h59 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_89 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_89 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_89 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_89 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_90 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h5a == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_90 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_90 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_90 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_90 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_91 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h5b == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_91 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_91 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_91 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_91 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_92 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h5c == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_92 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_92 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_92 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_92 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_93 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h5d == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_93 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_93 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_93 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_93 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_94 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h5e == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_94 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_94 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_94 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_94 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_95 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h5f == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_95 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_95 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_95 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_95 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_96 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h60 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_96 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_96 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_96 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_96 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_97 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h61 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_97 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_97 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_97 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_97 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_98 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h62 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_98 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_98 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_98 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_98 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_99 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h63 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_99 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_99 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_99 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_99 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_100 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h64 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_100 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_100 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_100 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_100 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_101 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h65 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_101 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_101 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_101 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_101 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_102 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h66 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_102 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_102 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_102 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_102 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_103 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h67 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_103 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_103 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_103 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_103 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_104 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h68 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_104 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_104 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_104 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_104 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_105 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h69 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_105 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_105 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_105 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_105 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_106 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h6a == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_106 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_106 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_106 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_106 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_107 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h6b == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_107 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_107 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_107 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_107 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_108 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h6c == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_108 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_108 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_108 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_108 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_109 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h6d == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_109 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_109 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_109 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_109 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_110 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h6e == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_110 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_110 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_110 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_110 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_111 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h6f == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_111 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_111 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_111 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_111 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_112 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h70 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_112 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_112 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_112 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_112 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_113 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h71 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_113 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_113 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_113 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_113 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_114 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h72 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_114 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_114 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_114 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_114 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_115 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h73 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_115 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_115 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_115 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_115 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_116 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h74 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_116 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_116 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_116 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_116 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_117 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h75 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_117 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_117 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_117 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_117 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_118 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h76 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_118 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_118 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_118 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_118 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_119 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h77 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_119 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_119 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_119 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_119 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_120 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h78 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_120 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_120 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_120 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_120 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_121 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h79 == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_121 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_121 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_121 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_121 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_122 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h7a == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_122 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_122 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_122 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_122 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_123 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h7b == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_123 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_123 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_123 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_123 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_124 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h7c == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_124 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_124 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_124 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_124 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_125 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h7d == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_125 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_125 <= tag_asid_regs_127;
      end else if (7'h7e == io_addr[10:4]) begin
        tag_asid_regs_125 <= tag_asid_regs_126;
      end else begin
        tag_asid_regs_125 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_126 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h7e == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_126 <= 8'h0;
      end else if (7'h7f == io_addr[10:4]) begin
        tag_asid_regs_126 <= tag_asid_regs_127;
      end else if (!(7'h7e == io_addr[10:4])) begin
        tag_asid_regs_126 <= _GEN_125;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[icache_tag.scala 33:34]
      tag_asid_regs_127 <= 8'h0; // @[icache_tag.scala 33:{40,40,40,40,40}]
    end else if (7'h7f == io_addr[10:4]) begin // @[icache_tag.scala 22:32]
      if (io_wen) begin
        tag_asid_regs_127 <= 8'h0;
      end else if (!(7'h7f == io_addr[10:4])) begin
        if (7'h7e == io_addr[10:4]) begin
          tag_asid_regs_127 <= tag_asid_regs_126;
        end else begin
          tag_asid_regs_127 <= _GEN_125;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tag_regs_0 = _RAND_0[21:0];
  _RAND_1 = {1{`RANDOM}};
  tag_regs_1 = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  tag_regs_2 = _RAND_2[21:0];
  _RAND_3 = {1{`RANDOM}};
  tag_regs_3 = _RAND_3[21:0];
  _RAND_4 = {1{`RANDOM}};
  tag_regs_4 = _RAND_4[21:0];
  _RAND_5 = {1{`RANDOM}};
  tag_regs_5 = _RAND_5[21:0];
  _RAND_6 = {1{`RANDOM}};
  tag_regs_6 = _RAND_6[21:0];
  _RAND_7 = {1{`RANDOM}};
  tag_regs_7 = _RAND_7[21:0];
  _RAND_8 = {1{`RANDOM}};
  tag_regs_8 = _RAND_8[21:0];
  _RAND_9 = {1{`RANDOM}};
  tag_regs_9 = _RAND_9[21:0];
  _RAND_10 = {1{`RANDOM}};
  tag_regs_10 = _RAND_10[21:0];
  _RAND_11 = {1{`RANDOM}};
  tag_regs_11 = _RAND_11[21:0];
  _RAND_12 = {1{`RANDOM}};
  tag_regs_12 = _RAND_12[21:0];
  _RAND_13 = {1{`RANDOM}};
  tag_regs_13 = _RAND_13[21:0];
  _RAND_14 = {1{`RANDOM}};
  tag_regs_14 = _RAND_14[21:0];
  _RAND_15 = {1{`RANDOM}};
  tag_regs_15 = _RAND_15[21:0];
  _RAND_16 = {1{`RANDOM}};
  tag_regs_16 = _RAND_16[21:0];
  _RAND_17 = {1{`RANDOM}};
  tag_regs_17 = _RAND_17[21:0];
  _RAND_18 = {1{`RANDOM}};
  tag_regs_18 = _RAND_18[21:0];
  _RAND_19 = {1{`RANDOM}};
  tag_regs_19 = _RAND_19[21:0];
  _RAND_20 = {1{`RANDOM}};
  tag_regs_20 = _RAND_20[21:0];
  _RAND_21 = {1{`RANDOM}};
  tag_regs_21 = _RAND_21[21:0];
  _RAND_22 = {1{`RANDOM}};
  tag_regs_22 = _RAND_22[21:0];
  _RAND_23 = {1{`RANDOM}};
  tag_regs_23 = _RAND_23[21:0];
  _RAND_24 = {1{`RANDOM}};
  tag_regs_24 = _RAND_24[21:0];
  _RAND_25 = {1{`RANDOM}};
  tag_regs_25 = _RAND_25[21:0];
  _RAND_26 = {1{`RANDOM}};
  tag_regs_26 = _RAND_26[21:0];
  _RAND_27 = {1{`RANDOM}};
  tag_regs_27 = _RAND_27[21:0];
  _RAND_28 = {1{`RANDOM}};
  tag_regs_28 = _RAND_28[21:0];
  _RAND_29 = {1{`RANDOM}};
  tag_regs_29 = _RAND_29[21:0];
  _RAND_30 = {1{`RANDOM}};
  tag_regs_30 = _RAND_30[21:0];
  _RAND_31 = {1{`RANDOM}};
  tag_regs_31 = _RAND_31[21:0];
  _RAND_32 = {1{`RANDOM}};
  tag_regs_32 = _RAND_32[21:0];
  _RAND_33 = {1{`RANDOM}};
  tag_regs_33 = _RAND_33[21:0];
  _RAND_34 = {1{`RANDOM}};
  tag_regs_34 = _RAND_34[21:0];
  _RAND_35 = {1{`RANDOM}};
  tag_regs_35 = _RAND_35[21:0];
  _RAND_36 = {1{`RANDOM}};
  tag_regs_36 = _RAND_36[21:0];
  _RAND_37 = {1{`RANDOM}};
  tag_regs_37 = _RAND_37[21:0];
  _RAND_38 = {1{`RANDOM}};
  tag_regs_38 = _RAND_38[21:0];
  _RAND_39 = {1{`RANDOM}};
  tag_regs_39 = _RAND_39[21:0];
  _RAND_40 = {1{`RANDOM}};
  tag_regs_40 = _RAND_40[21:0];
  _RAND_41 = {1{`RANDOM}};
  tag_regs_41 = _RAND_41[21:0];
  _RAND_42 = {1{`RANDOM}};
  tag_regs_42 = _RAND_42[21:0];
  _RAND_43 = {1{`RANDOM}};
  tag_regs_43 = _RAND_43[21:0];
  _RAND_44 = {1{`RANDOM}};
  tag_regs_44 = _RAND_44[21:0];
  _RAND_45 = {1{`RANDOM}};
  tag_regs_45 = _RAND_45[21:0];
  _RAND_46 = {1{`RANDOM}};
  tag_regs_46 = _RAND_46[21:0];
  _RAND_47 = {1{`RANDOM}};
  tag_regs_47 = _RAND_47[21:0];
  _RAND_48 = {1{`RANDOM}};
  tag_regs_48 = _RAND_48[21:0];
  _RAND_49 = {1{`RANDOM}};
  tag_regs_49 = _RAND_49[21:0];
  _RAND_50 = {1{`RANDOM}};
  tag_regs_50 = _RAND_50[21:0];
  _RAND_51 = {1{`RANDOM}};
  tag_regs_51 = _RAND_51[21:0];
  _RAND_52 = {1{`RANDOM}};
  tag_regs_52 = _RAND_52[21:0];
  _RAND_53 = {1{`RANDOM}};
  tag_regs_53 = _RAND_53[21:0];
  _RAND_54 = {1{`RANDOM}};
  tag_regs_54 = _RAND_54[21:0];
  _RAND_55 = {1{`RANDOM}};
  tag_regs_55 = _RAND_55[21:0];
  _RAND_56 = {1{`RANDOM}};
  tag_regs_56 = _RAND_56[21:0];
  _RAND_57 = {1{`RANDOM}};
  tag_regs_57 = _RAND_57[21:0];
  _RAND_58 = {1{`RANDOM}};
  tag_regs_58 = _RAND_58[21:0];
  _RAND_59 = {1{`RANDOM}};
  tag_regs_59 = _RAND_59[21:0];
  _RAND_60 = {1{`RANDOM}};
  tag_regs_60 = _RAND_60[21:0];
  _RAND_61 = {1{`RANDOM}};
  tag_regs_61 = _RAND_61[21:0];
  _RAND_62 = {1{`RANDOM}};
  tag_regs_62 = _RAND_62[21:0];
  _RAND_63 = {1{`RANDOM}};
  tag_regs_63 = _RAND_63[21:0];
  _RAND_64 = {1{`RANDOM}};
  tag_regs_64 = _RAND_64[21:0];
  _RAND_65 = {1{`RANDOM}};
  tag_regs_65 = _RAND_65[21:0];
  _RAND_66 = {1{`RANDOM}};
  tag_regs_66 = _RAND_66[21:0];
  _RAND_67 = {1{`RANDOM}};
  tag_regs_67 = _RAND_67[21:0];
  _RAND_68 = {1{`RANDOM}};
  tag_regs_68 = _RAND_68[21:0];
  _RAND_69 = {1{`RANDOM}};
  tag_regs_69 = _RAND_69[21:0];
  _RAND_70 = {1{`RANDOM}};
  tag_regs_70 = _RAND_70[21:0];
  _RAND_71 = {1{`RANDOM}};
  tag_regs_71 = _RAND_71[21:0];
  _RAND_72 = {1{`RANDOM}};
  tag_regs_72 = _RAND_72[21:0];
  _RAND_73 = {1{`RANDOM}};
  tag_regs_73 = _RAND_73[21:0];
  _RAND_74 = {1{`RANDOM}};
  tag_regs_74 = _RAND_74[21:0];
  _RAND_75 = {1{`RANDOM}};
  tag_regs_75 = _RAND_75[21:0];
  _RAND_76 = {1{`RANDOM}};
  tag_regs_76 = _RAND_76[21:0];
  _RAND_77 = {1{`RANDOM}};
  tag_regs_77 = _RAND_77[21:0];
  _RAND_78 = {1{`RANDOM}};
  tag_regs_78 = _RAND_78[21:0];
  _RAND_79 = {1{`RANDOM}};
  tag_regs_79 = _RAND_79[21:0];
  _RAND_80 = {1{`RANDOM}};
  tag_regs_80 = _RAND_80[21:0];
  _RAND_81 = {1{`RANDOM}};
  tag_regs_81 = _RAND_81[21:0];
  _RAND_82 = {1{`RANDOM}};
  tag_regs_82 = _RAND_82[21:0];
  _RAND_83 = {1{`RANDOM}};
  tag_regs_83 = _RAND_83[21:0];
  _RAND_84 = {1{`RANDOM}};
  tag_regs_84 = _RAND_84[21:0];
  _RAND_85 = {1{`RANDOM}};
  tag_regs_85 = _RAND_85[21:0];
  _RAND_86 = {1{`RANDOM}};
  tag_regs_86 = _RAND_86[21:0];
  _RAND_87 = {1{`RANDOM}};
  tag_regs_87 = _RAND_87[21:0];
  _RAND_88 = {1{`RANDOM}};
  tag_regs_88 = _RAND_88[21:0];
  _RAND_89 = {1{`RANDOM}};
  tag_regs_89 = _RAND_89[21:0];
  _RAND_90 = {1{`RANDOM}};
  tag_regs_90 = _RAND_90[21:0];
  _RAND_91 = {1{`RANDOM}};
  tag_regs_91 = _RAND_91[21:0];
  _RAND_92 = {1{`RANDOM}};
  tag_regs_92 = _RAND_92[21:0];
  _RAND_93 = {1{`RANDOM}};
  tag_regs_93 = _RAND_93[21:0];
  _RAND_94 = {1{`RANDOM}};
  tag_regs_94 = _RAND_94[21:0];
  _RAND_95 = {1{`RANDOM}};
  tag_regs_95 = _RAND_95[21:0];
  _RAND_96 = {1{`RANDOM}};
  tag_regs_96 = _RAND_96[21:0];
  _RAND_97 = {1{`RANDOM}};
  tag_regs_97 = _RAND_97[21:0];
  _RAND_98 = {1{`RANDOM}};
  tag_regs_98 = _RAND_98[21:0];
  _RAND_99 = {1{`RANDOM}};
  tag_regs_99 = _RAND_99[21:0];
  _RAND_100 = {1{`RANDOM}};
  tag_regs_100 = _RAND_100[21:0];
  _RAND_101 = {1{`RANDOM}};
  tag_regs_101 = _RAND_101[21:0];
  _RAND_102 = {1{`RANDOM}};
  tag_regs_102 = _RAND_102[21:0];
  _RAND_103 = {1{`RANDOM}};
  tag_regs_103 = _RAND_103[21:0];
  _RAND_104 = {1{`RANDOM}};
  tag_regs_104 = _RAND_104[21:0];
  _RAND_105 = {1{`RANDOM}};
  tag_regs_105 = _RAND_105[21:0];
  _RAND_106 = {1{`RANDOM}};
  tag_regs_106 = _RAND_106[21:0];
  _RAND_107 = {1{`RANDOM}};
  tag_regs_107 = _RAND_107[21:0];
  _RAND_108 = {1{`RANDOM}};
  tag_regs_108 = _RAND_108[21:0];
  _RAND_109 = {1{`RANDOM}};
  tag_regs_109 = _RAND_109[21:0];
  _RAND_110 = {1{`RANDOM}};
  tag_regs_110 = _RAND_110[21:0];
  _RAND_111 = {1{`RANDOM}};
  tag_regs_111 = _RAND_111[21:0];
  _RAND_112 = {1{`RANDOM}};
  tag_regs_112 = _RAND_112[21:0];
  _RAND_113 = {1{`RANDOM}};
  tag_regs_113 = _RAND_113[21:0];
  _RAND_114 = {1{`RANDOM}};
  tag_regs_114 = _RAND_114[21:0];
  _RAND_115 = {1{`RANDOM}};
  tag_regs_115 = _RAND_115[21:0];
  _RAND_116 = {1{`RANDOM}};
  tag_regs_116 = _RAND_116[21:0];
  _RAND_117 = {1{`RANDOM}};
  tag_regs_117 = _RAND_117[21:0];
  _RAND_118 = {1{`RANDOM}};
  tag_regs_118 = _RAND_118[21:0];
  _RAND_119 = {1{`RANDOM}};
  tag_regs_119 = _RAND_119[21:0];
  _RAND_120 = {1{`RANDOM}};
  tag_regs_120 = _RAND_120[21:0];
  _RAND_121 = {1{`RANDOM}};
  tag_regs_121 = _RAND_121[21:0];
  _RAND_122 = {1{`RANDOM}};
  tag_regs_122 = _RAND_122[21:0];
  _RAND_123 = {1{`RANDOM}};
  tag_regs_123 = _RAND_123[21:0];
  _RAND_124 = {1{`RANDOM}};
  tag_regs_124 = _RAND_124[21:0];
  _RAND_125 = {1{`RANDOM}};
  tag_regs_125 = _RAND_125[21:0];
  _RAND_126 = {1{`RANDOM}};
  tag_regs_126 = _RAND_126[21:0];
  _RAND_127 = {1{`RANDOM}};
  tag_regs_127 = _RAND_127[21:0];
  _RAND_128 = {1{`RANDOM}};
  tag_asid_regs_0 = _RAND_128[7:0];
  _RAND_129 = {1{`RANDOM}};
  tag_asid_regs_1 = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  tag_asid_regs_2 = _RAND_130[7:0];
  _RAND_131 = {1{`RANDOM}};
  tag_asid_regs_3 = _RAND_131[7:0];
  _RAND_132 = {1{`RANDOM}};
  tag_asid_regs_4 = _RAND_132[7:0];
  _RAND_133 = {1{`RANDOM}};
  tag_asid_regs_5 = _RAND_133[7:0];
  _RAND_134 = {1{`RANDOM}};
  tag_asid_regs_6 = _RAND_134[7:0];
  _RAND_135 = {1{`RANDOM}};
  tag_asid_regs_7 = _RAND_135[7:0];
  _RAND_136 = {1{`RANDOM}};
  tag_asid_regs_8 = _RAND_136[7:0];
  _RAND_137 = {1{`RANDOM}};
  tag_asid_regs_9 = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  tag_asid_regs_10 = _RAND_138[7:0];
  _RAND_139 = {1{`RANDOM}};
  tag_asid_regs_11 = _RAND_139[7:0];
  _RAND_140 = {1{`RANDOM}};
  tag_asid_regs_12 = _RAND_140[7:0];
  _RAND_141 = {1{`RANDOM}};
  tag_asid_regs_13 = _RAND_141[7:0];
  _RAND_142 = {1{`RANDOM}};
  tag_asid_regs_14 = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  tag_asid_regs_15 = _RAND_143[7:0];
  _RAND_144 = {1{`RANDOM}};
  tag_asid_regs_16 = _RAND_144[7:0];
  _RAND_145 = {1{`RANDOM}};
  tag_asid_regs_17 = _RAND_145[7:0];
  _RAND_146 = {1{`RANDOM}};
  tag_asid_regs_18 = _RAND_146[7:0];
  _RAND_147 = {1{`RANDOM}};
  tag_asid_regs_19 = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  tag_asid_regs_20 = _RAND_148[7:0];
  _RAND_149 = {1{`RANDOM}};
  tag_asid_regs_21 = _RAND_149[7:0];
  _RAND_150 = {1{`RANDOM}};
  tag_asid_regs_22 = _RAND_150[7:0];
  _RAND_151 = {1{`RANDOM}};
  tag_asid_regs_23 = _RAND_151[7:0];
  _RAND_152 = {1{`RANDOM}};
  tag_asid_regs_24 = _RAND_152[7:0];
  _RAND_153 = {1{`RANDOM}};
  tag_asid_regs_25 = _RAND_153[7:0];
  _RAND_154 = {1{`RANDOM}};
  tag_asid_regs_26 = _RAND_154[7:0];
  _RAND_155 = {1{`RANDOM}};
  tag_asid_regs_27 = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  tag_asid_regs_28 = _RAND_156[7:0];
  _RAND_157 = {1{`RANDOM}};
  tag_asid_regs_29 = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  tag_asid_regs_30 = _RAND_158[7:0];
  _RAND_159 = {1{`RANDOM}};
  tag_asid_regs_31 = _RAND_159[7:0];
  _RAND_160 = {1{`RANDOM}};
  tag_asid_regs_32 = _RAND_160[7:0];
  _RAND_161 = {1{`RANDOM}};
  tag_asid_regs_33 = _RAND_161[7:0];
  _RAND_162 = {1{`RANDOM}};
  tag_asid_regs_34 = _RAND_162[7:0];
  _RAND_163 = {1{`RANDOM}};
  tag_asid_regs_35 = _RAND_163[7:0];
  _RAND_164 = {1{`RANDOM}};
  tag_asid_regs_36 = _RAND_164[7:0];
  _RAND_165 = {1{`RANDOM}};
  tag_asid_regs_37 = _RAND_165[7:0];
  _RAND_166 = {1{`RANDOM}};
  tag_asid_regs_38 = _RAND_166[7:0];
  _RAND_167 = {1{`RANDOM}};
  tag_asid_regs_39 = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  tag_asid_regs_40 = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  tag_asid_regs_41 = _RAND_169[7:0];
  _RAND_170 = {1{`RANDOM}};
  tag_asid_regs_42 = _RAND_170[7:0];
  _RAND_171 = {1{`RANDOM}};
  tag_asid_regs_43 = _RAND_171[7:0];
  _RAND_172 = {1{`RANDOM}};
  tag_asid_regs_44 = _RAND_172[7:0];
  _RAND_173 = {1{`RANDOM}};
  tag_asid_regs_45 = _RAND_173[7:0];
  _RAND_174 = {1{`RANDOM}};
  tag_asid_regs_46 = _RAND_174[7:0];
  _RAND_175 = {1{`RANDOM}};
  tag_asid_regs_47 = _RAND_175[7:0];
  _RAND_176 = {1{`RANDOM}};
  tag_asid_regs_48 = _RAND_176[7:0];
  _RAND_177 = {1{`RANDOM}};
  tag_asid_regs_49 = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  tag_asid_regs_50 = _RAND_178[7:0];
  _RAND_179 = {1{`RANDOM}};
  tag_asid_regs_51 = _RAND_179[7:0];
  _RAND_180 = {1{`RANDOM}};
  tag_asid_regs_52 = _RAND_180[7:0];
  _RAND_181 = {1{`RANDOM}};
  tag_asid_regs_53 = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  tag_asid_regs_54 = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  tag_asid_regs_55 = _RAND_183[7:0];
  _RAND_184 = {1{`RANDOM}};
  tag_asid_regs_56 = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  tag_asid_regs_57 = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  tag_asid_regs_58 = _RAND_186[7:0];
  _RAND_187 = {1{`RANDOM}};
  tag_asid_regs_59 = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  tag_asid_regs_60 = _RAND_188[7:0];
  _RAND_189 = {1{`RANDOM}};
  tag_asid_regs_61 = _RAND_189[7:0];
  _RAND_190 = {1{`RANDOM}};
  tag_asid_regs_62 = _RAND_190[7:0];
  _RAND_191 = {1{`RANDOM}};
  tag_asid_regs_63 = _RAND_191[7:0];
  _RAND_192 = {1{`RANDOM}};
  tag_asid_regs_64 = _RAND_192[7:0];
  _RAND_193 = {1{`RANDOM}};
  tag_asid_regs_65 = _RAND_193[7:0];
  _RAND_194 = {1{`RANDOM}};
  tag_asid_regs_66 = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  tag_asid_regs_67 = _RAND_195[7:0];
  _RAND_196 = {1{`RANDOM}};
  tag_asid_regs_68 = _RAND_196[7:0];
  _RAND_197 = {1{`RANDOM}};
  tag_asid_regs_69 = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  tag_asid_regs_70 = _RAND_198[7:0];
  _RAND_199 = {1{`RANDOM}};
  tag_asid_regs_71 = _RAND_199[7:0];
  _RAND_200 = {1{`RANDOM}};
  tag_asid_regs_72 = _RAND_200[7:0];
  _RAND_201 = {1{`RANDOM}};
  tag_asid_regs_73 = _RAND_201[7:0];
  _RAND_202 = {1{`RANDOM}};
  tag_asid_regs_74 = _RAND_202[7:0];
  _RAND_203 = {1{`RANDOM}};
  tag_asid_regs_75 = _RAND_203[7:0];
  _RAND_204 = {1{`RANDOM}};
  tag_asid_regs_76 = _RAND_204[7:0];
  _RAND_205 = {1{`RANDOM}};
  tag_asid_regs_77 = _RAND_205[7:0];
  _RAND_206 = {1{`RANDOM}};
  tag_asid_regs_78 = _RAND_206[7:0];
  _RAND_207 = {1{`RANDOM}};
  tag_asid_regs_79 = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  tag_asid_regs_80 = _RAND_208[7:0];
  _RAND_209 = {1{`RANDOM}};
  tag_asid_regs_81 = _RAND_209[7:0];
  _RAND_210 = {1{`RANDOM}};
  tag_asid_regs_82 = _RAND_210[7:0];
  _RAND_211 = {1{`RANDOM}};
  tag_asid_regs_83 = _RAND_211[7:0];
  _RAND_212 = {1{`RANDOM}};
  tag_asid_regs_84 = _RAND_212[7:0];
  _RAND_213 = {1{`RANDOM}};
  tag_asid_regs_85 = _RAND_213[7:0];
  _RAND_214 = {1{`RANDOM}};
  tag_asid_regs_86 = _RAND_214[7:0];
  _RAND_215 = {1{`RANDOM}};
  tag_asid_regs_87 = _RAND_215[7:0];
  _RAND_216 = {1{`RANDOM}};
  tag_asid_regs_88 = _RAND_216[7:0];
  _RAND_217 = {1{`RANDOM}};
  tag_asid_regs_89 = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  tag_asid_regs_90 = _RAND_218[7:0];
  _RAND_219 = {1{`RANDOM}};
  tag_asid_regs_91 = _RAND_219[7:0];
  _RAND_220 = {1{`RANDOM}};
  tag_asid_regs_92 = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  tag_asid_regs_93 = _RAND_221[7:0];
  _RAND_222 = {1{`RANDOM}};
  tag_asid_regs_94 = _RAND_222[7:0];
  _RAND_223 = {1{`RANDOM}};
  tag_asid_regs_95 = _RAND_223[7:0];
  _RAND_224 = {1{`RANDOM}};
  tag_asid_regs_96 = _RAND_224[7:0];
  _RAND_225 = {1{`RANDOM}};
  tag_asid_regs_97 = _RAND_225[7:0];
  _RAND_226 = {1{`RANDOM}};
  tag_asid_regs_98 = _RAND_226[7:0];
  _RAND_227 = {1{`RANDOM}};
  tag_asid_regs_99 = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  tag_asid_regs_100 = _RAND_228[7:0];
  _RAND_229 = {1{`RANDOM}};
  tag_asid_regs_101 = _RAND_229[7:0];
  _RAND_230 = {1{`RANDOM}};
  tag_asid_regs_102 = _RAND_230[7:0];
  _RAND_231 = {1{`RANDOM}};
  tag_asid_regs_103 = _RAND_231[7:0];
  _RAND_232 = {1{`RANDOM}};
  tag_asid_regs_104 = _RAND_232[7:0];
  _RAND_233 = {1{`RANDOM}};
  tag_asid_regs_105 = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  tag_asid_regs_106 = _RAND_234[7:0];
  _RAND_235 = {1{`RANDOM}};
  tag_asid_regs_107 = _RAND_235[7:0];
  _RAND_236 = {1{`RANDOM}};
  tag_asid_regs_108 = _RAND_236[7:0];
  _RAND_237 = {1{`RANDOM}};
  tag_asid_regs_109 = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  tag_asid_regs_110 = _RAND_238[7:0];
  _RAND_239 = {1{`RANDOM}};
  tag_asid_regs_111 = _RAND_239[7:0];
  _RAND_240 = {1{`RANDOM}};
  tag_asid_regs_112 = _RAND_240[7:0];
  _RAND_241 = {1{`RANDOM}};
  tag_asid_regs_113 = _RAND_241[7:0];
  _RAND_242 = {1{`RANDOM}};
  tag_asid_regs_114 = _RAND_242[7:0];
  _RAND_243 = {1{`RANDOM}};
  tag_asid_regs_115 = _RAND_243[7:0];
  _RAND_244 = {1{`RANDOM}};
  tag_asid_regs_116 = _RAND_244[7:0];
  _RAND_245 = {1{`RANDOM}};
  tag_asid_regs_117 = _RAND_245[7:0];
  _RAND_246 = {1{`RANDOM}};
  tag_asid_regs_118 = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  tag_asid_regs_119 = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  tag_asid_regs_120 = _RAND_248[7:0];
  _RAND_249 = {1{`RANDOM}};
  tag_asid_regs_121 = _RAND_249[7:0];
  _RAND_250 = {1{`RANDOM}};
  tag_asid_regs_122 = _RAND_250[7:0];
  _RAND_251 = {1{`RANDOM}};
  tag_asid_regs_123 = _RAND_251[7:0];
  _RAND_252 = {1{`RANDOM}};
  tag_asid_regs_124 = _RAND_252[7:0];
  _RAND_253 = {1{`RANDOM}};
  tag_asid_regs_125 = _RAND_253[7:0];
  _RAND_254 = {1{`RANDOM}};
  tag_asid_regs_126 = _RAND_254[7:0];
  _RAND_255 = {1{`RANDOM}};
  tag_asid_regs_127 = _RAND_255[7:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    tag_regs_0 = 22'h0;
  end
  if (reset) begin
    tag_regs_1 = 22'h0;
  end
  if (reset) begin
    tag_regs_2 = 22'h0;
  end
  if (reset) begin
    tag_regs_3 = 22'h0;
  end
  if (reset) begin
    tag_regs_4 = 22'h0;
  end
  if (reset) begin
    tag_regs_5 = 22'h0;
  end
  if (reset) begin
    tag_regs_6 = 22'h0;
  end
  if (reset) begin
    tag_regs_7 = 22'h0;
  end
  if (reset) begin
    tag_regs_8 = 22'h0;
  end
  if (reset) begin
    tag_regs_9 = 22'h0;
  end
  if (reset) begin
    tag_regs_10 = 22'h0;
  end
  if (reset) begin
    tag_regs_11 = 22'h0;
  end
  if (reset) begin
    tag_regs_12 = 22'h0;
  end
  if (reset) begin
    tag_regs_13 = 22'h0;
  end
  if (reset) begin
    tag_regs_14 = 22'h0;
  end
  if (reset) begin
    tag_regs_15 = 22'h0;
  end
  if (reset) begin
    tag_regs_16 = 22'h0;
  end
  if (reset) begin
    tag_regs_17 = 22'h0;
  end
  if (reset) begin
    tag_regs_18 = 22'h0;
  end
  if (reset) begin
    tag_regs_19 = 22'h0;
  end
  if (reset) begin
    tag_regs_20 = 22'h0;
  end
  if (reset) begin
    tag_regs_21 = 22'h0;
  end
  if (reset) begin
    tag_regs_22 = 22'h0;
  end
  if (reset) begin
    tag_regs_23 = 22'h0;
  end
  if (reset) begin
    tag_regs_24 = 22'h0;
  end
  if (reset) begin
    tag_regs_25 = 22'h0;
  end
  if (reset) begin
    tag_regs_26 = 22'h0;
  end
  if (reset) begin
    tag_regs_27 = 22'h0;
  end
  if (reset) begin
    tag_regs_28 = 22'h0;
  end
  if (reset) begin
    tag_regs_29 = 22'h0;
  end
  if (reset) begin
    tag_regs_30 = 22'h0;
  end
  if (reset) begin
    tag_regs_31 = 22'h0;
  end
  if (reset) begin
    tag_regs_32 = 22'h0;
  end
  if (reset) begin
    tag_regs_33 = 22'h0;
  end
  if (reset) begin
    tag_regs_34 = 22'h0;
  end
  if (reset) begin
    tag_regs_35 = 22'h0;
  end
  if (reset) begin
    tag_regs_36 = 22'h0;
  end
  if (reset) begin
    tag_regs_37 = 22'h0;
  end
  if (reset) begin
    tag_regs_38 = 22'h0;
  end
  if (reset) begin
    tag_regs_39 = 22'h0;
  end
  if (reset) begin
    tag_regs_40 = 22'h0;
  end
  if (reset) begin
    tag_regs_41 = 22'h0;
  end
  if (reset) begin
    tag_regs_42 = 22'h0;
  end
  if (reset) begin
    tag_regs_43 = 22'h0;
  end
  if (reset) begin
    tag_regs_44 = 22'h0;
  end
  if (reset) begin
    tag_regs_45 = 22'h0;
  end
  if (reset) begin
    tag_regs_46 = 22'h0;
  end
  if (reset) begin
    tag_regs_47 = 22'h0;
  end
  if (reset) begin
    tag_regs_48 = 22'h0;
  end
  if (reset) begin
    tag_regs_49 = 22'h0;
  end
  if (reset) begin
    tag_regs_50 = 22'h0;
  end
  if (reset) begin
    tag_regs_51 = 22'h0;
  end
  if (reset) begin
    tag_regs_52 = 22'h0;
  end
  if (reset) begin
    tag_regs_53 = 22'h0;
  end
  if (reset) begin
    tag_regs_54 = 22'h0;
  end
  if (reset) begin
    tag_regs_55 = 22'h0;
  end
  if (reset) begin
    tag_regs_56 = 22'h0;
  end
  if (reset) begin
    tag_regs_57 = 22'h0;
  end
  if (reset) begin
    tag_regs_58 = 22'h0;
  end
  if (reset) begin
    tag_regs_59 = 22'h0;
  end
  if (reset) begin
    tag_regs_60 = 22'h0;
  end
  if (reset) begin
    tag_regs_61 = 22'h0;
  end
  if (reset) begin
    tag_regs_62 = 22'h0;
  end
  if (reset) begin
    tag_regs_63 = 22'h0;
  end
  if (reset) begin
    tag_regs_64 = 22'h0;
  end
  if (reset) begin
    tag_regs_65 = 22'h0;
  end
  if (reset) begin
    tag_regs_66 = 22'h0;
  end
  if (reset) begin
    tag_regs_67 = 22'h0;
  end
  if (reset) begin
    tag_regs_68 = 22'h0;
  end
  if (reset) begin
    tag_regs_69 = 22'h0;
  end
  if (reset) begin
    tag_regs_70 = 22'h0;
  end
  if (reset) begin
    tag_regs_71 = 22'h0;
  end
  if (reset) begin
    tag_regs_72 = 22'h0;
  end
  if (reset) begin
    tag_regs_73 = 22'h0;
  end
  if (reset) begin
    tag_regs_74 = 22'h0;
  end
  if (reset) begin
    tag_regs_75 = 22'h0;
  end
  if (reset) begin
    tag_regs_76 = 22'h0;
  end
  if (reset) begin
    tag_regs_77 = 22'h0;
  end
  if (reset) begin
    tag_regs_78 = 22'h0;
  end
  if (reset) begin
    tag_regs_79 = 22'h0;
  end
  if (reset) begin
    tag_regs_80 = 22'h0;
  end
  if (reset) begin
    tag_regs_81 = 22'h0;
  end
  if (reset) begin
    tag_regs_82 = 22'h0;
  end
  if (reset) begin
    tag_regs_83 = 22'h0;
  end
  if (reset) begin
    tag_regs_84 = 22'h0;
  end
  if (reset) begin
    tag_regs_85 = 22'h0;
  end
  if (reset) begin
    tag_regs_86 = 22'h0;
  end
  if (reset) begin
    tag_regs_87 = 22'h0;
  end
  if (reset) begin
    tag_regs_88 = 22'h0;
  end
  if (reset) begin
    tag_regs_89 = 22'h0;
  end
  if (reset) begin
    tag_regs_90 = 22'h0;
  end
  if (reset) begin
    tag_regs_91 = 22'h0;
  end
  if (reset) begin
    tag_regs_92 = 22'h0;
  end
  if (reset) begin
    tag_regs_93 = 22'h0;
  end
  if (reset) begin
    tag_regs_94 = 22'h0;
  end
  if (reset) begin
    tag_regs_95 = 22'h0;
  end
  if (reset) begin
    tag_regs_96 = 22'h0;
  end
  if (reset) begin
    tag_regs_97 = 22'h0;
  end
  if (reset) begin
    tag_regs_98 = 22'h0;
  end
  if (reset) begin
    tag_regs_99 = 22'h0;
  end
  if (reset) begin
    tag_regs_100 = 22'h0;
  end
  if (reset) begin
    tag_regs_101 = 22'h0;
  end
  if (reset) begin
    tag_regs_102 = 22'h0;
  end
  if (reset) begin
    tag_regs_103 = 22'h0;
  end
  if (reset) begin
    tag_regs_104 = 22'h0;
  end
  if (reset) begin
    tag_regs_105 = 22'h0;
  end
  if (reset) begin
    tag_regs_106 = 22'h0;
  end
  if (reset) begin
    tag_regs_107 = 22'h0;
  end
  if (reset) begin
    tag_regs_108 = 22'h0;
  end
  if (reset) begin
    tag_regs_109 = 22'h0;
  end
  if (reset) begin
    tag_regs_110 = 22'h0;
  end
  if (reset) begin
    tag_regs_111 = 22'h0;
  end
  if (reset) begin
    tag_regs_112 = 22'h0;
  end
  if (reset) begin
    tag_regs_113 = 22'h0;
  end
  if (reset) begin
    tag_regs_114 = 22'h0;
  end
  if (reset) begin
    tag_regs_115 = 22'h0;
  end
  if (reset) begin
    tag_regs_116 = 22'h0;
  end
  if (reset) begin
    tag_regs_117 = 22'h0;
  end
  if (reset) begin
    tag_regs_118 = 22'h0;
  end
  if (reset) begin
    tag_regs_119 = 22'h0;
  end
  if (reset) begin
    tag_regs_120 = 22'h0;
  end
  if (reset) begin
    tag_regs_121 = 22'h0;
  end
  if (reset) begin
    tag_regs_122 = 22'h0;
  end
  if (reset) begin
    tag_regs_123 = 22'h0;
  end
  if (reset) begin
    tag_regs_124 = 22'h0;
  end
  if (reset) begin
    tag_regs_125 = 22'h0;
  end
  if (reset) begin
    tag_regs_126 = 22'h0;
  end
  if (reset) begin
    tag_regs_127 = 22'h0;
  end
  if (reset) begin
    tag_asid_regs_0 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_1 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_2 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_3 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_4 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_5 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_6 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_7 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_8 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_9 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_10 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_11 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_12 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_13 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_14 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_15 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_16 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_17 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_18 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_19 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_20 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_21 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_22 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_23 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_24 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_25 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_26 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_27 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_28 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_29 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_30 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_31 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_32 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_33 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_34 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_35 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_36 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_37 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_38 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_39 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_40 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_41 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_42 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_43 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_44 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_45 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_46 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_47 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_48 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_49 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_50 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_51 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_52 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_53 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_54 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_55 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_56 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_57 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_58 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_59 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_60 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_61 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_62 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_63 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_64 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_65 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_66 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_67 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_68 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_69 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_70 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_71 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_72 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_73 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_74 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_75 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_76 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_77 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_78 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_79 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_80 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_81 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_82 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_83 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_84 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_85 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_86 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_87 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_88 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_89 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_90 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_91 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_92 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_93 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_94 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_95 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_96 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_97 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_98 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_99 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_100 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_101 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_102 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_103 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_104 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_105 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_106 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_107 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_108 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_109 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_110 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_111 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_112 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_113 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_114 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_115 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_116 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_117 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_118 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_119 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_120 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_121 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_122 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_123 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_124 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_125 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_126 = 8'h0;
  end
  if (reset) begin
    tag_asid_regs_127 = 8'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ysyx_sram_with_mask(
  input         clock,
  input  [7:0]  io_wea,
  input  [6:0]  io_addra,
  input  [63:0] io_dina,
  output [63:0] io_douta
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [127:0] S011HD1P_X32Y2D128_BW_Q; // @[ip_user.scala 140:22]
  wire  S011HD1P_X32Y2D128_BW_CLK; // @[ip_user.scala 140:22]
  wire  S011HD1P_X32Y2D128_BW_CEN; // @[ip_user.scala 140:22]
  wire  S011HD1P_X32Y2D128_BW_WEN; // @[ip_user.scala 140:22]
  wire [127:0] S011HD1P_X32Y2D128_BW_BWEN; // @[ip_user.scala 140:22]
  wire [5:0] S011HD1P_X32Y2D128_BW_A; // @[ip_user.scala 140:22]
  wire [127:0] S011HD1P_X32Y2D128_BW_D; // @[ip_user.scala 140:22]
  wire [127:0] final_write_data_1 = {io_dina, 64'h0}; // @[ip_user.scala 149:44]
  wire [7:0] ena_budle__0 = io_wea[0] ? 8'h0 : 8'hff; // @[ip_user.scala 154:35]
  wire [7:0] ena_budle__1 = io_wea[1] ? 8'h0 : 8'hff; // @[ip_user.scala 154:35]
  wire [7:0] ena_budle__2 = io_wea[2] ? 8'h0 : 8'hff; // @[ip_user.scala 154:35]
  wire [7:0] ena_budle__3 = io_wea[3] ? 8'h0 : 8'hff; // @[ip_user.scala 154:35]
  wire [7:0] ena_budle__4 = io_wea[4] ? 8'h0 : 8'hff; // @[ip_user.scala 154:35]
  wire [7:0] ena_budle__5 = io_wea[5] ? 8'h0 : 8'hff; // @[ip_user.scala 154:35]
  wire [7:0] ena_budle__6 = io_wea[6] ? 8'h0 : 8'hff; // @[ip_user.scala 154:35]
  wire [7:0] ena_budle__7 = io_wea[7] ? 8'h0 : 8'hff; // @[ip_user.scala 154:35]
  wire [63:0] _final_ena_data_0_T_2 = {ena_budle__7,ena_budle__6,ena_budle__5,ena_budle__4,ena_budle__3,ena_budle__2,
    ena_budle__1,ena_budle__0}; // @[ip_user.scala 156:96]
  wire [63:0] final_ena_data_0 = ~io_addra[0] ? _final_ena_data_0_T_2 : 64'hffffffffffffffff; // @[ip_user.scala 156:38]
  wire [63:0] final_ena_data_1 = io_addra[0] ? _final_ena_data_0_T_2 : 64'hffffffffffffffff; // @[ip_user.scala 156:38]
  wire [127:0] final_write_data_0 = {{64'd0}, io_dina}; // @[ip_user.scala 146:32 149:33]
  reg [6:0] addr_reg; // @[ip_user.scala 164:28]
  wire  shift_num = addr_reg[0]; // @[ip_user.scala 165:30]
  wire [63:0] sram_data_bundle_0 = S011HD1P_X32Y2D128_BW_Q[63:0]; // @[ip_user.scala 168:42]
  wire [63:0] sram_data_bundle_1 = S011HD1P_X32Y2D128_BW_Q[127:64]; // @[ip_user.scala 168:42]
  S011HD1P_X32Y2D128_BW S011HD1P_X32Y2D128_BW ( // @[ip_user.scala 140:22]
    .Q(S011HD1P_X32Y2D128_BW_Q),
    .CLK(S011HD1P_X32Y2D128_BW_CLK),
    .CEN(S011HD1P_X32Y2D128_BW_CEN),
    .WEN(S011HD1P_X32Y2D128_BW_WEN),
    .BWEN(S011HD1P_X32Y2D128_BW_BWEN),
    .A(S011HD1P_X32Y2D128_BW_A),
    .D(S011HD1P_X32Y2D128_BW_D)
  );
  assign io_douta = shift_num ? sram_data_bundle_1 : sram_data_bundle_0; // @[ip_user.scala 170:{14,14}]
  assign S011HD1P_X32Y2D128_BW_CLK = clock; // @[ip_user.scala 142:23]
  assign S011HD1P_X32Y2D128_BW_CEN = 1'h0; // @[ip_user.scala 141:17]
  assign S011HD1P_X32Y2D128_BW_WEN = io_wea == 8'h0; // @[ip_user.scala 143:24]
  assign S011HD1P_X32Y2D128_BW_BWEN = {final_ena_data_1,final_ena_data_0}; // @[ip_user.scala 162:33]
  assign S011HD1P_X32Y2D128_BW_A = io_addra[6:1]; // @[ip_user.scala 163:23]
  assign S011HD1P_X32Y2D128_BW_D = io_addra[0] ? final_write_data_1 : final_write_data_0; // @[ip_user.scala 161:{12,12}]
  always @(posedge clock) begin
    addr_reg <= io_addra; // @[ip_user.scala 164:28]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr_reg = _RAND_0[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module icache_data(
  input         clock,
  input  [7:0]  io_wen,
  input  [63:0] io_addr,
  input  [63:0] io_wdata,
  output [39:0] io_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  icache_data_ram_0_clock; // @[icache_data.scala 31:35]
  wire [7:0] icache_data_ram_0_io_wea; // @[icache_data.scala 31:35]
  wire [6:0] icache_data_ram_0_io_addra; // @[icache_data.scala 31:35]
  wire [63:0] icache_data_ram_0_io_dina; // @[icache_data.scala 31:35]
  wire [63:0] icache_data_ram_0_io_douta; // @[icache_data.scala 31:35]
  reg [63:0] addr_reg; // @[icache_data.scala 36:27]
  wire [31:0] get_data = addr_reg[2] ? icache_data_ram_0_io_douta[63:32] : icache_data_ram_0_io_douta[31:0]; // @[icache_data.scala 38:26]
  wire [6:0] io_rdata_opD = get_data[6:0]; // @[macros.scala 524:24]
  wire [2:0] io_rdata_Funct3D = get_data[14:12]; // @[macros.scala 525:28]
  wire [1:0] _io_rdata_T_3 = 3'h1 == io_rdata_Funct3D ? 2'h2 : {{1'd0}, 3'h0 == io_rdata_Funct3D}; // @[Mux.scala 81:58]
  wire [2:0] _io_rdata_T_5 = 3'h4 == io_rdata_Funct3D ? 3'h4 : {{1'd0}, _io_rdata_T_3}; // @[Mux.scala 81:58]
  wire [3:0] _io_rdata_T_7 = 3'h5 == io_rdata_Funct3D ? 4'h8 : {{1'd0}, _io_rdata_T_5}; // @[Mux.scala 81:58]
  wire [4:0] _io_rdata_T_9 = 3'h6 == io_rdata_Funct3D ? 5'h10 : {{1'd0}, _io_rdata_T_7}; // @[Mux.scala 81:58]
  wire [5:0] _io_rdata_T_11 = 3'h7 == io_rdata_Funct3D ? 6'h20 : {{1'd0}, _io_rdata_T_9}; // @[Mux.scala 81:58]
  wire [5:0] _io_rdata_T_13 = 7'h63 == io_rdata_opD ? _io_rdata_T_11 : 6'h0; // @[Mux.scala 81:58]
  wire  _io_rdata_T_16 = io_rdata_opD == 7'h67 & io_rdata_Funct3D == 3'h0; // @[macros.scala 497:30]
  wire  _io_rdata_T_18 = _io_rdata_T_16 | io_rdata_opD == 7'h6f; // @[macros.scala 502:27]
  wire  _io_rdata_T_19 = io_rdata_opD == 7'h63; // @[macros.scala 520:13]
  wire [32:0] io_rdata_lo = {_io_rdata_T_19,get_data}; // @[Cat.scala 31:58]
  wire [6:0] io_rdata_hi = {_io_rdata_T_13,_io_rdata_T_18}; // @[Cat.scala 31:58]
  ysyx_sram_with_mask icache_data_ram_0 ( // @[icache_data.scala 31:35]
    .clock(icache_data_ram_0_clock),
    .io_wea(icache_data_ram_0_io_wea),
    .io_addra(icache_data_ram_0_io_addra),
    .io_dina(icache_data_ram_0_io_dina),
    .io_douta(icache_data_ram_0_io_douta)
  );
  assign io_rdata = {io_rdata_hi,io_rdata_lo}; // @[Cat.scala 31:58]
  assign icache_data_ram_0_clock = clock;
  assign icache_data_ram_0_io_wea = io_wen; // @[icache_data.scala 33:31]
  assign icache_data_ram_0_io_addra = io_addr[10:4]; // @[icache_data.scala 34:42]
  assign icache_data_ram_0_io_dina = io_wdata; // @[icache_data.scala 35:31]
  always @(posedge clock) begin
    addr_reg <= io_addr; // @[icache_data.scala 36:27]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  addr_reg = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module inst_cache(
  input         clock,
  input         reset,
  output [63:0] io_port_araddr,
  output [3:0]  io_port_arlen,
  output [1:0]  io_port_arburst,
  output        io_port_arvalid,
  input         io_port_arready,
  input  [63:0] io_port_rdata,
  input         io_port_rlast,
  input         io_port_rvalid,
  input         io_stage2_flush,
  output        io_stage2_stall,
  input         io_stage1_valid_flush,
  input         io_inst_ready_to_use,
  input         io_inst_buffer_full,
  output [63:0] io_v_addr_for_tlb,
  input  [63:0] io_p_addr_for_tlb,
  input         io_sram_req,
  input  [63:0] io_sram_addr,
  output [1:0]  io_sram_write_en,
  output [39:0] io_sram_rdata_L,
  input         io_sram_cache,
  input         io_tag_valid_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [63:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [63:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [63:0] _RAND_142;
`endif // RANDOMIZE_REG_INIT
  wire  icache_tag_clock; // @[inst_cache.scala 81:34]
  wire  icache_tag_reset; // @[inst_cache.scala 81:34]
  wire  icache_tag_io_wen; // @[inst_cache.scala 81:34]
  wire [20:0] icache_tag_io_wdata; // @[inst_cache.scala 81:34]
  wire [63:0] icache_tag_io_addr; // @[inst_cache.scala 81:34]
  wire  icache_tag_io_hit; // @[inst_cache.scala 81:34]
  wire  icache_tag_io_valid; // @[inst_cache.scala 81:34]
  wire  icache_tag_io_tag_all_flush; // @[inst_cache.scala 81:34]
  wire  icache_tag_1_clock; // @[inst_cache.scala 83:34]
  wire  icache_tag_1_reset; // @[inst_cache.scala 83:34]
  wire  icache_tag_1_io_wen; // @[inst_cache.scala 83:34]
  wire [20:0] icache_tag_1_io_wdata; // @[inst_cache.scala 83:34]
  wire [63:0] icache_tag_1_io_addr; // @[inst_cache.scala 83:34]
  wire  icache_tag_1_io_hit; // @[inst_cache.scala 83:34]
  wire  icache_tag_1_io_valid; // @[inst_cache.scala 83:34]
  wire  icache_tag_1_io_tag_all_flush; // @[inst_cache.scala 83:34]
  wire  icache_data_clock; // @[inst_cache.scala 89:55]
  wire [7:0] icache_data_io_wen; // @[inst_cache.scala 89:55]
  wire [63:0] icache_data_io_addr; // @[inst_cache.scala 89:55]
  wire [63:0] icache_data_io_wdata; // @[inst_cache.scala 89:55]
  wire [39:0] icache_data_io_rdata; // @[inst_cache.scala 89:55]
  wire  icache_data_1_clock; // @[inst_cache.scala 89:55]
  wire [7:0] icache_data_1_io_wen; // @[inst_cache.scala 89:55]
  wire [63:0] icache_data_1_io_addr; // @[inst_cache.scala 89:55]
  wire [63:0] icache_data_1_io_wdata; // @[inst_cache.scala 89:55]
  wire [39:0] icache_data_1_io_rdata; // @[inst_cache.scala 89:55]
  wire  icache_data_2_clock; // @[inst_cache.scala 90:55]
  wire [7:0] icache_data_2_io_wen; // @[inst_cache.scala 90:55]
  wire [63:0] icache_data_2_io_addr; // @[inst_cache.scala 90:55]
  wire [63:0] icache_data_2_io_wdata; // @[inst_cache.scala 90:55]
  wire [39:0] icache_data_2_io_rdata; // @[inst_cache.scala 90:55]
  wire  icache_data_3_clock; // @[inst_cache.scala 90:55]
  wire [7:0] icache_data_3_io_wen; // @[inst_cache.scala 90:55]
  wire [63:0] icache_data_3_io_addr; // @[inst_cache.scala 90:55]
  wire [63:0] icache_data_3_io_wdata; // @[inst_cache.scala 90:55]
  wire [39:0] icache_data_3_io_rdata; // @[inst_cache.scala 90:55]
  reg  lru_0; // @[inst_cache.scala 74:22]
  reg  lru_1; // @[inst_cache.scala 74:22]
  reg  lru_2; // @[inst_cache.scala 74:22]
  reg  lru_3; // @[inst_cache.scala 74:22]
  reg  lru_4; // @[inst_cache.scala 74:22]
  reg  lru_5; // @[inst_cache.scala 74:22]
  reg  lru_6; // @[inst_cache.scala 74:22]
  reg  lru_7; // @[inst_cache.scala 74:22]
  reg  lru_8; // @[inst_cache.scala 74:22]
  reg  lru_9; // @[inst_cache.scala 74:22]
  reg  lru_10; // @[inst_cache.scala 74:22]
  reg  lru_11; // @[inst_cache.scala 74:22]
  reg  lru_12; // @[inst_cache.scala 74:22]
  reg  lru_13; // @[inst_cache.scala 74:22]
  reg  lru_14; // @[inst_cache.scala 74:22]
  reg  lru_15; // @[inst_cache.scala 74:22]
  reg  lru_16; // @[inst_cache.scala 74:22]
  reg  lru_17; // @[inst_cache.scala 74:22]
  reg  lru_18; // @[inst_cache.scala 74:22]
  reg  lru_19; // @[inst_cache.scala 74:22]
  reg  lru_20; // @[inst_cache.scala 74:22]
  reg  lru_21; // @[inst_cache.scala 74:22]
  reg  lru_22; // @[inst_cache.scala 74:22]
  reg  lru_23; // @[inst_cache.scala 74:22]
  reg  lru_24; // @[inst_cache.scala 74:22]
  reg  lru_25; // @[inst_cache.scala 74:22]
  reg  lru_26; // @[inst_cache.scala 74:22]
  reg  lru_27; // @[inst_cache.scala 74:22]
  reg  lru_28; // @[inst_cache.scala 74:22]
  reg  lru_29; // @[inst_cache.scala 74:22]
  reg  lru_30; // @[inst_cache.scala 74:22]
  reg  lru_31; // @[inst_cache.scala 74:22]
  reg  lru_32; // @[inst_cache.scala 74:22]
  reg  lru_33; // @[inst_cache.scala 74:22]
  reg  lru_34; // @[inst_cache.scala 74:22]
  reg  lru_35; // @[inst_cache.scala 74:22]
  reg  lru_36; // @[inst_cache.scala 74:22]
  reg  lru_37; // @[inst_cache.scala 74:22]
  reg  lru_38; // @[inst_cache.scala 74:22]
  reg  lru_39; // @[inst_cache.scala 74:22]
  reg  lru_40; // @[inst_cache.scala 74:22]
  reg  lru_41; // @[inst_cache.scala 74:22]
  reg  lru_42; // @[inst_cache.scala 74:22]
  reg  lru_43; // @[inst_cache.scala 74:22]
  reg  lru_44; // @[inst_cache.scala 74:22]
  reg  lru_45; // @[inst_cache.scala 74:22]
  reg  lru_46; // @[inst_cache.scala 74:22]
  reg  lru_47; // @[inst_cache.scala 74:22]
  reg  lru_48; // @[inst_cache.scala 74:22]
  reg  lru_49; // @[inst_cache.scala 74:22]
  reg  lru_50; // @[inst_cache.scala 74:22]
  reg  lru_51; // @[inst_cache.scala 74:22]
  reg  lru_52; // @[inst_cache.scala 74:22]
  reg  lru_53; // @[inst_cache.scala 74:22]
  reg  lru_54; // @[inst_cache.scala 74:22]
  reg  lru_55; // @[inst_cache.scala 74:22]
  reg  lru_56; // @[inst_cache.scala 74:22]
  reg  lru_57; // @[inst_cache.scala 74:22]
  reg  lru_58; // @[inst_cache.scala 74:22]
  reg  lru_59; // @[inst_cache.scala 74:22]
  reg  lru_60; // @[inst_cache.scala 74:22]
  reg  lru_61; // @[inst_cache.scala 74:22]
  reg  lru_62; // @[inst_cache.scala 74:22]
  reg  lru_63; // @[inst_cache.scala 74:22]
  reg  lru_64; // @[inst_cache.scala 74:22]
  reg  lru_65; // @[inst_cache.scala 74:22]
  reg  lru_66; // @[inst_cache.scala 74:22]
  reg  lru_67; // @[inst_cache.scala 74:22]
  reg  lru_68; // @[inst_cache.scala 74:22]
  reg  lru_69; // @[inst_cache.scala 74:22]
  reg  lru_70; // @[inst_cache.scala 74:22]
  reg  lru_71; // @[inst_cache.scala 74:22]
  reg  lru_72; // @[inst_cache.scala 74:22]
  reg  lru_73; // @[inst_cache.scala 74:22]
  reg  lru_74; // @[inst_cache.scala 74:22]
  reg  lru_75; // @[inst_cache.scala 74:22]
  reg  lru_76; // @[inst_cache.scala 74:22]
  reg  lru_77; // @[inst_cache.scala 74:22]
  reg  lru_78; // @[inst_cache.scala 74:22]
  reg  lru_79; // @[inst_cache.scala 74:22]
  reg  lru_80; // @[inst_cache.scala 74:22]
  reg  lru_81; // @[inst_cache.scala 74:22]
  reg  lru_82; // @[inst_cache.scala 74:22]
  reg  lru_83; // @[inst_cache.scala 74:22]
  reg  lru_84; // @[inst_cache.scala 74:22]
  reg  lru_85; // @[inst_cache.scala 74:22]
  reg  lru_86; // @[inst_cache.scala 74:22]
  reg  lru_87; // @[inst_cache.scala 74:22]
  reg  lru_88; // @[inst_cache.scala 74:22]
  reg  lru_89; // @[inst_cache.scala 74:22]
  reg  lru_90; // @[inst_cache.scala 74:22]
  reg  lru_91; // @[inst_cache.scala 74:22]
  reg  lru_92; // @[inst_cache.scala 74:22]
  reg  lru_93; // @[inst_cache.scala 74:22]
  reg  lru_94; // @[inst_cache.scala 74:22]
  reg  lru_95; // @[inst_cache.scala 74:22]
  reg  lru_96; // @[inst_cache.scala 74:22]
  reg  lru_97; // @[inst_cache.scala 74:22]
  reg  lru_98; // @[inst_cache.scala 74:22]
  reg  lru_99; // @[inst_cache.scala 74:22]
  reg  lru_100; // @[inst_cache.scala 74:22]
  reg  lru_101; // @[inst_cache.scala 74:22]
  reg  lru_102; // @[inst_cache.scala 74:22]
  reg  lru_103; // @[inst_cache.scala 74:22]
  reg  lru_104; // @[inst_cache.scala 74:22]
  reg  lru_105; // @[inst_cache.scala 74:22]
  reg  lru_106; // @[inst_cache.scala 74:22]
  reg  lru_107; // @[inst_cache.scala 74:22]
  reg  lru_108; // @[inst_cache.scala 74:22]
  reg  lru_109; // @[inst_cache.scala 74:22]
  reg  lru_110; // @[inst_cache.scala 74:22]
  reg  lru_111; // @[inst_cache.scala 74:22]
  reg  lru_112; // @[inst_cache.scala 74:22]
  reg  lru_113; // @[inst_cache.scala 74:22]
  reg  lru_114; // @[inst_cache.scala 74:22]
  reg  lru_115; // @[inst_cache.scala 74:22]
  reg  lru_116; // @[inst_cache.scala 74:22]
  reg  lru_117; // @[inst_cache.scala 74:22]
  reg  lru_118; // @[inst_cache.scala 74:22]
  reg  lru_119; // @[inst_cache.scala 74:22]
  reg  lru_120; // @[inst_cache.scala 74:22]
  reg  lru_121; // @[inst_cache.scala 74:22]
  reg  lru_122; // @[inst_cache.scala 74:22]
  reg  lru_123; // @[inst_cache.scala 74:22]
  reg  lru_124; // @[inst_cache.scala 74:22]
  reg  lru_125; // @[inst_cache.scala 74:22]
  reg  lru_126; // @[inst_cache.scala 74:22]
  reg  lru_127; // @[inst_cache.scala 74:22]
  reg [3:0] work_state; // @[inst_cache.scala 101:29]
  reg [2:0] write_counter; // @[inst_cache.scala 103:33]
  reg [39:0] wait_data_L; // @[inst_cache.scala 104:31]
  wire  stage1_flush = ~io_sram_req & io_stage1_valid_flush; // @[inst_cache.scala 108:35]
  reg  stage1_stall_reg; // @[inst_cache.scala 115:35]
  reg [63:0] stage1_addr_line_mapping; // @[Reg.scala 28:20]
  reg [63:0] stage1_sram_phy_addr_reg; // @[inst_cache.scala 119:43]
  reg  stage1_sram_cache_reg; // @[Reg.scala 28:20]
  wire  _stage1_sram_req_reg_T_1 = io_sram_req | stage1_flush; // @[inst_cache.scala 121:106]
  reg  stage1_sram_req_reg; // @[Reg.scala 28:20]
  reg  stage1_finished; // @[inst_cache.scala 124:34]
  wire  _stage1_finished_T_1 = work_state == 4'h7; // @[inst_cache.scala 140:67]
  wire  _stage1_finished_T_2 = work_state == 4'h3; // @[inst_cache.scala 140:103]
  wire  _access_work_state_T = work_state == 4'h2; // @[inst_cache.scala 244:41]
  wire  _access_work_state_T_6 = io_port_rlast & io_port_rvalid; // @[inst_cache.scala 245:71]
  wire [2:0] _access_work_state_T_7 = io_port_rlast & io_port_rvalid ? 3'h4 : 3'h3; // @[inst_cache.scala 245:49]
  wire  _access_work_state_T_8 = work_state == 4'h4; // @[inst_cache.scala 246:23]
  wire  _hit_T = icache_tag_io_hit; // @[inst_cache.scala 171:33]
  wire  _hit_T_2 = icache_tag_io_hit & icache_tag_io_valid; // @[inst_cache.scala 171:40]
  wire  _hit_T_3 = icache_tag_1_io_hit; // @[inst_cache.scala 172:27]
  wire  _hit_T_5 = icache_tag_1_io_hit & icache_tag_1_io_valid; // @[inst_cache.scala 172:34]
  wire  hit = icache_tag_io_hit & icache_tag_io_valid | _hit_T_5; // @[inst_cache.scala 171:70]
  wire [2:0] _access_work_state_T_13 = stage1_finished ? 3'h4 : 3'h2; // @[inst_cache.scala 246:145]
  wire [2:0] _access_work_state_T_14 = stage1_sram_cache_reg ? 3'h1 : _access_work_state_T_13; // @[inst_cache.scala 246:99]
  wire [2:0] _access_work_state_T_15 = stage1_sram_req_reg ? _access_work_state_T_14 : 3'h1; // @[inst_cache.scala 246:68]
  wire [2:0] _access_work_state_T_18 = stage1_finished ? 3'h4 : 3'h5; // @[inst_cache.scala 247:79]
  wire [2:0] _access_work_state_T_20 = stage1_sram_cache_reg ? _access_work_state_T_18 : _access_work_state_T_13; // @[inst_cache.scala 247:46]
  wire [2:0] _access_work_state_T_21 = stage1_sram_req_reg ? _access_work_state_T_20 : 3'h1; // @[inst_cache.scala 247:15]
  wire [2:0] _access_work_state_T_22 = hit ? _access_work_state_T_15 : _access_work_state_T_21; // @[inst_cache.scala 246:46]
  wire  _access_work_state_T_23 = work_state == 4'h1; // @[inst_cache.scala 249:23]
  wire [1:0] _access_work_state_T_28 = stage1_sram_cache_reg ? 2'h1 : 2'h2; // @[inst_cache.scala 249:95]
  wire [1:0] _access_work_state_T_29 = stage1_sram_req_reg ? _access_work_state_T_28 : 2'h1; // @[inst_cache.scala 249:64]
  wire [2:0] _access_work_state_T_32 = stage1_sram_cache_reg ? 3'h5 : 3'h2; // @[inst_cache.scala 250:46]
  wire [2:0] _access_work_state_T_33 = stage1_sram_req_reg ? _access_work_state_T_32 : 3'h1; // @[inst_cache.scala 250:15]
  wire [2:0] _access_work_state_T_34 = hit ? {{1'd0}, _access_work_state_T_29} : _access_work_state_T_33; // @[inst_cache.scala 249:42]
  wire  _access_work_state_T_35 = work_state == 4'h5; // @[inst_cache.scala 251:23]
  wire  _access_work_state_T_38 = work_state == 4'h6; // @[inst_cache.scala 252:23]
  wire [3:0] _access_work_state_T_42 = _access_work_state_T_6 ? 4'h7 : work_state; // @[inst_cache.scala 252:54]
  wire [3:0] _access_work_state_T_44 = _stage1_finished_T_1 ? 4'h4 : work_state; // @[inst_cache.scala 253:12]
  wire [3:0] _access_work_state_T_45 = work_state == 4'h6 ? _access_work_state_T_42 : _access_work_state_T_44; // @[inst_cache.scala 252:12]
  wire [3:0] _access_work_state_T_46 = work_state == 4'h5 & io_port_arready ? 4'h6 : _access_work_state_T_45; // @[inst_cache.scala 251:12]
  wire [3:0] _access_work_state_T_47 = work_state == 4'h1 ? {{1'd0}, _access_work_state_T_34} : _access_work_state_T_46; // @[inst_cache.scala 249:12]
  wire [3:0] _access_work_state_T_48 = work_state == 4'h4 ? {{1'd0}, _access_work_state_T_22} : _access_work_state_T_47; // @[inst_cache.scala 246:12]
  wire [3:0] _access_work_state_T_49 = _stage1_finished_T_2 ? {{1'd0}, _access_work_state_T_7} : _access_work_state_T_48
    ; // @[inst_cache.scala 245:12]
  wire [3:0] access_work_state = work_state == 4'h2 & io_port_arready ? 4'h3 : _access_work_state_T_49; // @[inst_cache.scala 244:30]
  wire  _stage2_stall_T = access_work_state == 4'h1; // @[inst_cache.scala 145:40]
  wire  _stage2_stall_T_5 = ~io_inst_buffer_full; // @[inst_cache.scala 146:11]
  wire  stage2_stall = (access_work_state == 4'h1 | access_work_state == 4'h4) & _stage2_stall_T_5; // @[inst_cache.scala 145:129]
  wire [6:0] decoder_inst_data_0_opD = io_port_rdata[6:0]; // @[macros.scala 524:24]
  wire [2:0] decoder_inst_data_0_Funct3D = io_port_rdata[14:12]; // @[macros.scala 525:28]
  wire [1:0] _decoder_inst_data_0_T_4 = 3'h1 == decoder_inst_data_0_Funct3D ? 2'h2 : {{1'd0}, 3'h0 ==
    decoder_inst_data_0_Funct3D}; // @[Mux.scala 81:58]
  wire [2:0] _decoder_inst_data_0_T_6 = 3'h4 == decoder_inst_data_0_Funct3D ? 3'h4 : {{1'd0}, _decoder_inst_data_0_T_4}; // @[Mux.scala 81:58]
  wire [3:0] _decoder_inst_data_0_T_8 = 3'h5 == decoder_inst_data_0_Funct3D ? 4'h8 : {{1'd0}, _decoder_inst_data_0_T_6}; // @[Mux.scala 81:58]
  wire [4:0] _decoder_inst_data_0_T_10 = 3'h6 == decoder_inst_data_0_Funct3D ? 5'h10 : {{1'd0}, _decoder_inst_data_0_T_8
    }; // @[Mux.scala 81:58]
  wire [5:0] _decoder_inst_data_0_T_12 = 3'h7 == decoder_inst_data_0_Funct3D ? 6'h20 : {{1'd0},
    _decoder_inst_data_0_T_10}; // @[Mux.scala 81:58]
  wire [5:0] _decoder_inst_data_0_T_14 = 7'h63 == decoder_inst_data_0_opD ? _decoder_inst_data_0_T_12 : 6'h0; // @[Mux.scala 81:58]
  wire  _decoder_inst_data_0_T_18 = decoder_inst_data_0_opD == 7'h67 & decoder_inst_data_0_Funct3D == 3'h0; // @[macros.scala 497:30]
  wire  _decoder_inst_data_0_T_20 = _decoder_inst_data_0_T_18 | decoder_inst_data_0_opD == 7'h6f; // @[macros.scala 502:27]
  wire  _decoder_inst_data_0_T_22 = decoder_inst_data_0_opD == 7'h63; // @[macros.scala 520:13]
  wire [39:0] decoder_inst_data_0 = {_decoder_inst_data_0_T_14,_decoder_inst_data_0_T_20,_decoder_inst_data_0_T_22,
    io_port_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [6:0] decoder_inst_data_1_opD = io_port_rdata[38:32]; // @[macros.scala 524:24]
  wire [2:0] decoder_inst_data_1_Funct3D = io_port_rdata[46:44]; // @[macros.scala 525:28]
  wire [1:0] _decoder_inst_data_1_T_4 = 3'h1 == decoder_inst_data_1_Funct3D ? 2'h2 : {{1'd0}, 3'h0 ==
    decoder_inst_data_1_Funct3D}; // @[Mux.scala 81:58]
  wire [2:0] _decoder_inst_data_1_T_6 = 3'h4 == decoder_inst_data_1_Funct3D ? 3'h4 : {{1'd0}, _decoder_inst_data_1_T_4}; // @[Mux.scala 81:58]
  wire [3:0] _decoder_inst_data_1_T_8 = 3'h5 == decoder_inst_data_1_Funct3D ? 4'h8 : {{1'd0}, _decoder_inst_data_1_T_6}; // @[Mux.scala 81:58]
  wire [4:0] _decoder_inst_data_1_T_10 = 3'h6 == decoder_inst_data_1_Funct3D ? 5'h10 : {{1'd0}, _decoder_inst_data_1_T_8
    }; // @[Mux.scala 81:58]
  wire [5:0] _decoder_inst_data_1_T_12 = 3'h7 == decoder_inst_data_1_Funct3D ? 6'h20 : {{1'd0},
    _decoder_inst_data_1_T_10}; // @[Mux.scala 81:58]
  wire [5:0] _decoder_inst_data_1_T_14 = 7'h63 == decoder_inst_data_1_opD ? _decoder_inst_data_1_T_12 : 6'h0; // @[Mux.scala 81:58]
  wire  _decoder_inst_data_1_T_18 = decoder_inst_data_1_opD == 7'h67 & decoder_inst_data_1_Funct3D == 3'h0; // @[macros.scala 497:30]
  wire  _decoder_inst_data_1_T_20 = _decoder_inst_data_1_T_18 | decoder_inst_data_1_opD == 7'h6f; // @[macros.scala 502:27]
  wire  _decoder_inst_data_1_T_22 = decoder_inst_data_1_opD == 7'h63; // @[macros.scala 520:13]
  wire [39:0] decoder_inst_data_1 = {_decoder_inst_data_1_T_14,_decoder_inst_data_1_T_20,_decoder_inst_data_1_T_22,
    io_port_rdata[63:32]}; // @[Cat.scala 31:58]
  wire [39:0] decoder_inst_data = stage1_addr_line_mapping[2] ? decoder_inst_data_1 : decoder_inst_data_0; // @[inst_cache.scala 156:33]
  wire  _GEN_4 = 7'h1 == stage1_addr_line_mapping[10:4] ? lru_1 : lru_0; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_5 = 7'h2 == stage1_addr_line_mapping[10:4] ? lru_2 : _GEN_4; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_6 = 7'h3 == stage1_addr_line_mapping[10:4] ? lru_3 : _GEN_5; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_7 = 7'h4 == stage1_addr_line_mapping[10:4] ? lru_4 : _GEN_6; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_8 = 7'h5 == stage1_addr_line_mapping[10:4] ? lru_5 : _GEN_7; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_9 = 7'h6 == stage1_addr_line_mapping[10:4] ? lru_6 : _GEN_8; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_10 = 7'h7 == stage1_addr_line_mapping[10:4] ? lru_7 : _GEN_9; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_11 = 7'h8 == stage1_addr_line_mapping[10:4] ? lru_8 : _GEN_10; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_12 = 7'h9 == stage1_addr_line_mapping[10:4] ? lru_9 : _GEN_11; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_13 = 7'ha == stage1_addr_line_mapping[10:4] ? lru_10 : _GEN_12; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_14 = 7'hb == stage1_addr_line_mapping[10:4] ? lru_11 : _GEN_13; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_15 = 7'hc == stage1_addr_line_mapping[10:4] ? lru_12 : _GEN_14; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_16 = 7'hd == stage1_addr_line_mapping[10:4] ? lru_13 : _GEN_15; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_17 = 7'he == stage1_addr_line_mapping[10:4] ? lru_14 : _GEN_16; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_18 = 7'hf == stage1_addr_line_mapping[10:4] ? lru_15 : _GEN_17; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_19 = 7'h10 == stage1_addr_line_mapping[10:4] ? lru_16 : _GEN_18; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_20 = 7'h11 == stage1_addr_line_mapping[10:4] ? lru_17 : _GEN_19; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_21 = 7'h12 == stage1_addr_line_mapping[10:4] ? lru_18 : _GEN_20; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_22 = 7'h13 == stage1_addr_line_mapping[10:4] ? lru_19 : _GEN_21; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_23 = 7'h14 == stage1_addr_line_mapping[10:4] ? lru_20 : _GEN_22; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_24 = 7'h15 == stage1_addr_line_mapping[10:4] ? lru_21 : _GEN_23; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_25 = 7'h16 == stage1_addr_line_mapping[10:4] ? lru_22 : _GEN_24; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_26 = 7'h17 == stage1_addr_line_mapping[10:4] ? lru_23 : _GEN_25; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_27 = 7'h18 == stage1_addr_line_mapping[10:4] ? lru_24 : _GEN_26; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_28 = 7'h19 == stage1_addr_line_mapping[10:4] ? lru_25 : _GEN_27; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_29 = 7'h1a == stage1_addr_line_mapping[10:4] ? lru_26 : _GEN_28; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_30 = 7'h1b == stage1_addr_line_mapping[10:4] ? lru_27 : _GEN_29; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_31 = 7'h1c == stage1_addr_line_mapping[10:4] ? lru_28 : _GEN_30; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_32 = 7'h1d == stage1_addr_line_mapping[10:4] ? lru_29 : _GEN_31; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_33 = 7'h1e == stage1_addr_line_mapping[10:4] ? lru_30 : _GEN_32; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_34 = 7'h1f == stage1_addr_line_mapping[10:4] ? lru_31 : _GEN_33; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_35 = 7'h20 == stage1_addr_line_mapping[10:4] ? lru_32 : _GEN_34; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_36 = 7'h21 == stage1_addr_line_mapping[10:4] ? lru_33 : _GEN_35; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_37 = 7'h22 == stage1_addr_line_mapping[10:4] ? lru_34 : _GEN_36; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_38 = 7'h23 == stage1_addr_line_mapping[10:4] ? lru_35 : _GEN_37; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_39 = 7'h24 == stage1_addr_line_mapping[10:4] ? lru_36 : _GEN_38; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_40 = 7'h25 == stage1_addr_line_mapping[10:4] ? lru_37 : _GEN_39; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_41 = 7'h26 == stage1_addr_line_mapping[10:4] ? lru_38 : _GEN_40; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_42 = 7'h27 == stage1_addr_line_mapping[10:4] ? lru_39 : _GEN_41; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_43 = 7'h28 == stage1_addr_line_mapping[10:4] ? lru_40 : _GEN_42; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_44 = 7'h29 == stage1_addr_line_mapping[10:4] ? lru_41 : _GEN_43; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_45 = 7'h2a == stage1_addr_line_mapping[10:4] ? lru_42 : _GEN_44; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_46 = 7'h2b == stage1_addr_line_mapping[10:4] ? lru_43 : _GEN_45; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_47 = 7'h2c == stage1_addr_line_mapping[10:4] ? lru_44 : _GEN_46; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_48 = 7'h2d == stage1_addr_line_mapping[10:4] ? lru_45 : _GEN_47; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_49 = 7'h2e == stage1_addr_line_mapping[10:4] ? lru_46 : _GEN_48; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_50 = 7'h2f == stage1_addr_line_mapping[10:4] ? lru_47 : _GEN_49; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_51 = 7'h30 == stage1_addr_line_mapping[10:4] ? lru_48 : _GEN_50; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_52 = 7'h31 == stage1_addr_line_mapping[10:4] ? lru_49 : _GEN_51; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_53 = 7'h32 == stage1_addr_line_mapping[10:4] ? lru_50 : _GEN_52; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_54 = 7'h33 == stage1_addr_line_mapping[10:4] ? lru_51 : _GEN_53; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_55 = 7'h34 == stage1_addr_line_mapping[10:4] ? lru_52 : _GEN_54; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_56 = 7'h35 == stage1_addr_line_mapping[10:4] ? lru_53 : _GEN_55; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_57 = 7'h36 == stage1_addr_line_mapping[10:4] ? lru_54 : _GEN_56; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_58 = 7'h37 == stage1_addr_line_mapping[10:4] ? lru_55 : _GEN_57; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_59 = 7'h38 == stage1_addr_line_mapping[10:4] ? lru_56 : _GEN_58; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_60 = 7'h39 == stage1_addr_line_mapping[10:4] ? lru_57 : _GEN_59; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_61 = 7'h3a == stage1_addr_line_mapping[10:4] ? lru_58 : _GEN_60; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_62 = 7'h3b == stage1_addr_line_mapping[10:4] ? lru_59 : _GEN_61; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_63 = 7'h3c == stage1_addr_line_mapping[10:4] ? lru_60 : _GEN_62; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_64 = 7'h3d == stage1_addr_line_mapping[10:4] ? lru_61 : _GEN_63; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_65 = 7'h3e == stage1_addr_line_mapping[10:4] ? lru_62 : _GEN_64; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_66 = 7'h3f == stage1_addr_line_mapping[10:4] ? lru_63 : _GEN_65; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_67 = 7'h40 == stage1_addr_line_mapping[10:4] ? lru_64 : _GEN_66; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_68 = 7'h41 == stage1_addr_line_mapping[10:4] ? lru_65 : _GEN_67; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_69 = 7'h42 == stage1_addr_line_mapping[10:4] ? lru_66 : _GEN_68; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_70 = 7'h43 == stage1_addr_line_mapping[10:4] ? lru_67 : _GEN_69; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_71 = 7'h44 == stage1_addr_line_mapping[10:4] ? lru_68 : _GEN_70; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_72 = 7'h45 == stage1_addr_line_mapping[10:4] ? lru_69 : _GEN_71; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_73 = 7'h46 == stage1_addr_line_mapping[10:4] ? lru_70 : _GEN_72; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_74 = 7'h47 == stage1_addr_line_mapping[10:4] ? lru_71 : _GEN_73; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_75 = 7'h48 == stage1_addr_line_mapping[10:4] ? lru_72 : _GEN_74; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_76 = 7'h49 == stage1_addr_line_mapping[10:4] ? lru_73 : _GEN_75; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_77 = 7'h4a == stage1_addr_line_mapping[10:4] ? lru_74 : _GEN_76; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_78 = 7'h4b == stage1_addr_line_mapping[10:4] ? lru_75 : _GEN_77; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_79 = 7'h4c == stage1_addr_line_mapping[10:4] ? lru_76 : _GEN_78; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_80 = 7'h4d == stage1_addr_line_mapping[10:4] ? lru_77 : _GEN_79; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_81 = 7'h4e == stage1_addr_line_mapping[10:4] ? lru_78 : _GEN_80; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_82 = 7'h4f == stage1_addr_line_mapping[10:4] ? lru_79 : _GEN_81; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_83 = 7'h50 == stage1_addr_line_mapping[10:4] ? lru_80 : _GEN_82; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_84 = 7'h51 == stage1_addr_line_mapping[10:4] ? lru_81 : _GEN_83; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_85 = 7'h52 == stage1_addr_line_mapping[10:4] ? lru_82 : _GEN_84; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_86 = 7'h53 == stage1_addr_line_mapping[10:4] ? lru_83 : _GEN_85; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_87 = 7'h54 == stage1_addr_line_mapping[10:4] ? lru_84 : _GEN_86; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_88 = 7'h55 == stage1_addr_line_mapping[10:4] ? lru_85 : _GEN_87; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_89 = 7'h56 == stage1_addr_line_mapping[10:4] ? lru_86 : _GEN_88; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_90 = 7'h57 == stage1_addr_line_mapping[10:4] ? lru_87 : _GEN_89; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_91 = 7'h58 == stage1_addr_line_mapping[10:4] ? lru_88 : _GEN_90; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_92 = 7'h59 == stage1_addr_line_mapping[10:4] ? lru_89 : _GEN_91; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_93 = 7'h5a == stage1_addr_line_mapping[10:4] ? lru_90 : _GEN_92; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_94 = 7'h5b == stage1_addr_line_mapping[10:4] ? lru_91 : _GEN_93; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_95 = 7'h5c == stage1_addr_line_mapping[10:4] ? lru_92 : _GEN_94; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_96 = 7'h5d == stage1_addr_line_mapping[10:4] ? lru_93 : _GEN_95; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_97 = 7'h5e == stage1_addr_line_mapping[10:4] ? lru_94 : _GEN_96; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_98 = 7'h5f == stage1_addr_line_mapping[10:4] ? lru_95 : _GEN_97; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_99 = 7'h60 == stage1_addr_line_mapping[10:4] ? lru_96 : _GEN_98; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_100 = 7'h61 == stage1_addr_line_mapping[10:4] ? lru_97 : _GEN_99; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_101 = 7'h62 == stage1_addr_line_mapping[10:4] ? lru_98 : _GEN_100; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_102 = 7'h63 == stage1_addr_line_mapping[10:4] ? lru_99 : _GEN_101; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_103 = 7'h64 == stage1_addr_line_mapping[10:4] ? lru_100 : _GEN_102; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_104 = 7'h65 == stage1_addr_line_mapping[10:4] ? lru_101 : _GEN_103; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_105 = 7'h66 == stage1_addr_line_mapping[10:4] ? lru_102 : _GEN_104; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_106 = 7'h67 == stage1_addr_line_mapping[10:4] ? lru_103 : _GEN_105; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_107 = 7'h68 == stage1_addr_line_mapping[10:4] ? lru_104 : _GEN_106; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_108 = 7'h69 == stage1_addr_line_mapping[10:4] ? lru_105 : _GEN_107; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_109 = 7'h6a == stage1_addr_line_mapping[10:4] ? lru_106 : _GEN_108; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_110 = 7'h6b == stage1_addr_line_mapping[10:4] ? lru_107 : _GEN_109; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_111 = 7'h6c == stage1_addr_line_mapping[10:4] ? lru_108 : _GEN_110; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_112 = 7'h6d == stage1_addr_line_mapping[10:4] ? lru_109 : _GEN_111; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_113 = 7'h6e == stage1_addr_line_mapping[10:4] ? lru_110 : _GEN_112; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_114 = 7'h6f == stage1_addr_line_mapping[10:4] ? lru_111 : _GEN_113; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_115 = 7'h70 == stage1_addr_line_mapping[10:4] ? lru_112 : _GEN_114; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_116 = 7'h71 == stage1_addr_line_mapping[10:4] ? lru_113 : _GEN_115; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_117 = 7'h72 == stage1_addr_line_mapping[10:4] ? lru_114 : _GEN_116; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_118 = 7'h73 == stage1_addr_line_mapping[10:4] ? lru_115 : _GEN_117; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_119 = 7'h74 == stage1_addr_line_mapping[10:4] ? lru_116 : _GEN_118; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_120 = 7'h75 == stage1_addr_line_mapping[10:4] ? lru_117 : _GEN_119; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_121 = 7'h76 == stage1_addr_line_mapping[10:4] ? lru_118 : _GEN_120; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_122 = 7'h77 == stage1_addr_line_mapping[10:4] ? lru_119 : _GEN_121; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_123 = 7'h78 == stage1_addr_line_mapping[10:4] ? lru_120 : _GEN_122; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_124 = 7'h79 == stage1_addr_line_mapping[10:4] ? lru_121 : _GEN_123; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_125 = 7'h7a == stage1_addr_line_mapping[10:4] ? lru_122 : _GEN_124; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_126 = 7'h7b == stage1_addr_line_mapping[10:4] ? lru_123 : _GEN_125; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_127 = 7'h7c == stage1_addr_line_mapping[10:4] ? lru_124 : _GEN_126; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_128 = 7'h7d == stage1_addr_line_mapping[10:4] ? lru_125 : _GEN_127; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_129 = 7'h7e == stage1_addr_line_mapping[10:4] ? lru_126 : _GEN_128; // @[inst_cache.scala 176:{12,12}]
  wire  _GEN_130 = 7'h7f == stage1_addr_line_mapping[10:4] ? lru_127 : _GEN_129; // @[inst_cache.scala 176:{12,12}]
  wire  _lru_T_4 = _hit_T_3 ? 1'h0 : _GEN_130; // @[inst_cache.scala 176:12]
  wire  _lru_T_5 = _hit_T | _lru_T_4; // @[inst_cache.scala 175:12]
  wire  _lru_T_8 = ~_GEN_130; // @[inst_cache.scala 177:46]
  reg [63:0] stage2_sram_addr_reg; // @[inst_cache.scala 182:39]
  reg  stage2_sram_req_reg; // @[inst_cache.scala 189:38]
  reg  stage2_hit0_reg; // @[inst_cache.scala 193:34]
  reg [1:0] stage2_write_en_reg; // @[inst_cache.scala 210:38]
  wire [39:0] icache_data_way0_0_rdata = icache_data_io_rdata; // @[inst_cache.scala 89:{36,36}]
  wire [39:0] icache_data_way0_1_rdata = icache_data_1_io_rdata; // @[inst_cache.scala 89:{36,36}]
  wire [39:0] _GEN_516 = stage2_sram_addr_reg[3] ? icache_data_way0_1_rdata : icache_data_way0_0_rdata; // @[inst_cache.scala 221:{25,25}]
  wire [39:0] icache_data_way1_0_rdata = icache_data_2_io_rdata; // @[inst_cache.scala 90:{36,36}]
  wire [39:0] icache_data_way1_1_rdata = icache_data_3_io_rdata; // @[inst_cache.scala 90:{36,36}]
  wire [39:0] _GEN_518 = stage2_sram_addr_reg[3] ? icache_data_way1_1_rdata : icache_data_way1_0_rdata; // @[inst_cache.scala 221:{25,25}]
  wire [39:0] hit_word_L = stage2_hit0_reg ? _GEN_516 : _GEN_518; // @[inst_cache.scala 221:25]
  reg  has_stage2_stall; // @[inst_cache.scala 223:35]
  reg [39:0] sram_rdata_L_Reg; // @[inst_cache.scala 226:35]
  wire [39:0] _access_sram_rdata_L_T_2 = _access_work_state_T_23 ? hit_word_L : 40'h0; // @[inst_cache.scala 229:84]
  wire [39:0] access_sram_rdata_L = _access_work_state_T_8 ? wait_data_L : _access_sram_rdata_L_T_2; // @[inst_cache.scala 229:35]
  wire  _icache_data_way0_0_wen_T_2 = _access_work_state_T_38 & io_port_rvalid; // @[inst_cache.scala 236:119]
  wire  _icache_data_way0_0_wen_T_6 = write_counter == 3'h0; // @[inst_cache.scala 237:69]
  wire  _icache_data_way0_0_wen_T_7 = _icache_data_way0_0_wen_T_2 & _lru_T_8 & write_counter == 3'h0; // @[inst_cache.scala 237:52]
  wire  _icache_data_way0_1_wen_T_6 = write_counter == 3'h1; // @[inst_cache.scala 237:69]
  wire  _icache_data_way0_1_wen_T_7 = _icache_data_way0_0_wen_T_2 & _lru_T_8 & write_counter == 3'h1; // @[inst_cache.scala 237:52]
  wire  _icache_data_way1_0_wen_T_7 = _icache_data_way0_0_wen_T_2 & _GEN_130 & _icache_data_way0_0_wen_T_6; // @[inst_cache.scala 239:52]
  wire  _icache_data_way1_1_wen_T_7 = _icache_data_way0_0_wen_T_2 & _GEN_130 & _icache_data_way0_1_wen_T_6; // @[inst_cache.scala 239:52]
  wire [2:0] _GEN_1287 = {{2'd0}, stage1_addr_line_mapping[3]}; // @[inst_cache.scala 259:95]
  wire [2:0] _write_counter_T_8 = write_counter + 3'h1; // @[inst_cache.scala 264:196]
  wire [21:0] _T_13 = {1'h1,stage1_addr_line_mapping[31:11]}; // @[Cat.scala 31:58]
  wire [21:0] _T_14 = _stage1_finished_T_1 ? _T_13 : 22'h0; // @[inst_cache.scala 267:30]
  wire [63:0] _io_port_araddr_T_3 = {stage1_sram_phy_addr_reg[63:4],4'h0}; // @[Cat.scala 31:58]
  wire [63:0] _io_port_araddr_T_4 = _access_work_state_T_35 ? _io_port_araddr_T_3 : 64'h0; // @[inst_cache.scala 278:12]
  wire  _io_sram_write_en_T_3 = ~stage2_sram_req_reg & stage2_sram_addr_reg[1:0] != 2'h0; // @[inst_cache.scala 317:31]
  wire [1:0] _io_sram_write_en_T_5 = stage2_sram_req_reg | _io_sram_write_en_T_3 ? stage2_write_en_reg : 2'h0; // @[inst_cache.scala 316:57]
  icache_tag icache_tag ( // @[inst_cache.scala 81:34]
    .clock(icache_tag_clock),
    .reset(icache_tag_reset),
    .io_wen(icache_tag_io_wen),
    .io_wdata(icache_tag_io_wdata),
    .io_addr(icache_tag_io_addr),
    .io_hit(icache_tag_io_hit),
    .io_valid(icache_tag_io_valid),
    .io_tag_all_flush(icache_tag_io_tag_all_flush)
  );
  icache_tag icache_tag_1 ( // @[inst_cache.scala 83:34]
    .clock(icache_tag_1_clock),
    .reset(icache_tag_1_reset),
    .io_wen(icache_tag_1_io_wen),
    .io_wdata(icache_tag_1_io_wdata),
    .io_addr(icache_tag_1_io_addr),
    .io_hit(icache_tag_1_io_hit),
    .io_valid(icache_tag_1_io_valid),
    .io_tag_all_flush(icache_tag_1_io_tag_all_flush)
  );
  icache_data icache_data ( // @[inst_cache.scala 89:55]
    .clock(icache_data_clock),
    .io_wen(icache_data_io_wen),
    .io_addr(icache_data_io_addr),
    .io_wdata(icache_data_io_wdata),
    .io_rdata(icache_data_io_rdata)
  );
  icache_data icache_data_1 ( // @[inst_cache.scala 89:55]
    .clock(icache_data_1_clock),
    .io_wen(icache_data_1_io_wen),
    .io_addr(icache_data_1_io_addr),
    .io_wdata(icache_data_1_io_wdata),
    .io_rdata(icache_data_1_io_rdata)
  );
  icache_data icache_data_2 ( // @[inst_cache.scala 90:55]
    .clock(icache_data_2_clock),
    .io_wen(icache_data_2_io_wen),
    .io_addr(icache_data_2_io_addr),
    .io_wdata(icache_data_2_io_wdata),
    .io_rdata(icache_data_2_io_rdata)
  );
  icache_data icache_data_3 ( // @[inst_cache.scala 90:55]
    .clock(icache_data_3_clock),
    .io_wen(icache_data_3_io_wen),
    .io_addr(icache_data_3_io_addr),
    .io_wdata(icache_data_3_io_wdata),
    .io_rdata(icache_data_3_io_rdata)
  );
  assign io_port_araddr = _access_work_state_T ? stage1_sram_phy_addr_reg : _io_port_araddr_T_4; // @[inst_cache.scala 277:26]
  assign io_port_arlen = {{3'd0}, stage1_sram_cache_reg}; // @[inst_cache.scala 280:20]
  assign io_port_arburst = {{1'd0}, stage1_sram_cache_reg}; // @[inst_cache.scala 282:21]
  assign io_port_arvalid = _access_work_state_T | _access_work_state_T_35; // @[inst_cache.scala 287:59]
  assign io_stage2_stall = (access_work_state == 4'h1 | access_work_state == 4'h4) & _stage2_stall_T_5; // @[inst_cache.scala 145:129]
  assign io_v_addr_for_tlb = stage1_addr_line_mapping; // @[inst_cache.scala 134:23]
  assign io_sram_write_en = io_inst_buffer_full ? 2'h0 : _io_sram_write_en_T_5; // @[inst_cache.scala 316:28]
  assign io_sram_rdata_L = _stage2_stall_T_5 & has_stage2_stall ? access_sram_rdata_L : sram_rdata_L_Reg; // @[inst_cache.scala 241:27]
  assign icache_tag_clock = clock;
  assign icache_tag_reset = reset;
  assign icache_tag_io_wen = _stage1_finished_T_1 & _lru_T_8; // @[inst_cache.scala 265:63]
  assign icache_tag_io_wdata = _T_14[20:0]; // @[inst_cache.scala 267:24]
  assign icache_tag_io_addr = stage1_addr_line_mapping; // @[inst_cache.scala 151:25]
  assign icache_tag_io_tag_all_flush = io_tag_valid_flush; // @[inst_cache.scala 87:32]
  assign icache_tag_1_clock = clock;
  assign icache_tag_1_reset = reset;
  assign icache_tag_1_io_wen = _stage1_finished_T_1 & _GEN_130; // @[inst_cache.scala 266:63]
  assign icache_tag_1_io_wdata = _T_14[20:0]; // @[inst_cache.scala 268:24]
  assign icache_tag_1_io_addr = stage1_addr_line_mapping; // @[inst_cache.scala 152:25]
  assign icache_tag_1_io_tag_all_flush = io_tag_valid_flush; // @[inst_cache.scala 88:32]
  assign icache_data_clock = clock;
  assign icache_data_io_wen = _icache_data_way0_0_wen_T_7 ? 8'hff : 8'h0; // @[inst_cache.scala 236:79]
  assign icache_data_io_addr = stage1_addr_line_mapping; // @[inst_cache.scala 161:34 89:36]
  assign icache_data_io_wdata = {io_port_rdata[63:32],io_port_rdata[31:0]}; // @[Cat.scala 31:58]
  assign icache_data_1_clock = clock;
  assign icache_data_1_io_wen = _icache_data_way0_1_wen_T_7 ? 8'hff : 8'h0; // @[inst_cache.scala 236:79]
  assign icache_data_1_io_addr = stage1_addr_line_mapping; // @[inst_cache.scala 161:34 89:36]
  assign icache_data_1_io_wdata = {io_port_rdata[63:32],io_port_rdata[31:0]}; // @[Cat.scala 31:58]
  assign icache_data_2_clock = clock;
  assign icache_data_2_io_wen = _icache_data_way1_0_wen_T_7 ? 8'hff : 8'h0; // @[inst_cache.scala 238:79]
  assign icache_data_2_io_addr = stage1_addr_line_mapping; // @[inst_cache.scala 166:34 90:36]
  assign icache_data_2_io_wdata = {io_port_rdata[63:32],io_port_rdata[31:0]}; // @[Cat.scala 31:58]
  assign icache_data_3_clock = clock;
  assign icache_data_3_io_wen = _icache_data_way1_1_wen_T_7 ? 8'hff : 8'h0; // @[inst_cache.scala 238:79]
  assign icache_data_3_io_addr = stage1_addr_line_mapping; // @[inst_cache.scala 166:34 90:36]
  assign icache_data_3_io_wdata = {io_port_rdata[63:32],io_port_rdata[31:0]}; // @[Cat.scala 31:58]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_0 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h0 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_0 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_0 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_0 <= lru_127;
      end else begin
        lru_0 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_1 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h1 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_1 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_1 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_1 <= lru_127;
      end else begin
        lru_1 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_2 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h2 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_2 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_2 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_2 <= lru_127;
      end else begin
        lru_2 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_3 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h3 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_3 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_3 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_3 <= lru_127;
      end else begin
        lru_3 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_4 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h4 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_4 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_4 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_4 <= lru_127;
      end else begin
        lru_4 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_5 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h5 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_5 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_5 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_5 <= lru_127;
      end else begin
        lru_5 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_6 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h6 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_6 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_6 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_6 <= lru_127;
      end else begin
        lru_6 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_7 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h7 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_7 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_7 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_7 <= lru_127;
      end else begin
        lru_7 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_8 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h8 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_8 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_8 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_8 <= lru_127;
      end else begin
        lru_8 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_9 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h9 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_9 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_9 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_9 <= lru_127;
      end else begin
        lru_9 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_10 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'ha == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_10 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_10 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_10 <= lru_127;
      end else begin
        lru_10 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_11 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'hb == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_11 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_11 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_11 <= lru_127;
      end else begin
        lru_11 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_12 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'hc == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_12 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_12 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_12 <= lru_127;
      end else begin
        lru_12 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_13 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'hd == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_13 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_13 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_13 <= lru_127;
      end else begin
        lru_13 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_14 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'he == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_14 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_14 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_14 <= lru_127;
      end else begin
        lru_14 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_15 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'hf == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_15 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_15 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_15 <= lru_127;
      end else begin
        lru_15 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_16 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h10 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_16 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_16 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_16 <= lru_127;
      end else begin
        lru_16 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_17 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h11 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_17 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_17 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_17 <= lru_127;
      end else begin
        lru_17 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_18 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h12 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_18 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_18 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_18 <= lru_127;
      end else begin
        lru_18 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_19 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h13 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_19 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_19 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_19 <= lru_127;
      end else begin
        lru_19 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_20 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h14 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_20 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_20 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_20 <= lru_127;
      end else begin
        lru_20 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_21 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h15 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_21 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_21 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_21 <= lru_127;
      end else begin
        lru_21 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_22 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h16 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_22 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_22 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_22 <= lru_127;
      end else begin
        lru_22 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_23 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h17 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_23 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_23 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_23 <= lru_127;
      end else begin
        lru_23 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_24 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h18 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_24 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_24 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_24 <= lru_127;
      end else begin
        lru_24 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_25 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h19 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_25 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_25 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_25 <= lru_127;
      end else begin
        lru_25 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_26 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h1a == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_26 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_26 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_26 <= lru_127;
      end else begin
        lru_26 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_27 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h1b == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_27 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_27 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_27 <= lru_127;
      end else begin
        lru_27 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_28 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h1c == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_28 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_28 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_28 <= lru_127;
      end else begin
        lru_28 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_29 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h1d == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_29 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_29 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_29 <= lru_127;
      end else begin
        lru_29 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_30 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h1e == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_30 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_30 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_30 <= lru_127;
      end else begin
        lru_30 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_31 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h1f == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_31 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_31 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_31 <= lru_127;
      end else begin
        lru_31 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_32 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h20 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_32 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_32 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_32 <= lru_127;
      end else begin
        lru_32 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_33 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h21 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_33 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_33 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_33 <= lru_127;
      end else begin
        lru_33 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_34 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h22 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_34 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_34 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_34 <= lru_127;
      end else begin
        lru_34 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_35 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h23 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_35 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_35 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_35 <= lru_127;
      end else begin
        lru_35 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_36 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h24 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_36 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_36 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_36 <= lru_127;
      end else begin
        lru_36 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_37 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h25 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_37 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_37 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_37 <= lru_127;
      end else begin
        lru_37 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_38 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h26 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_38 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_38 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_38 <= lru_127;
      end else begin
        lru_38 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_39 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h27 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_39 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_39 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_39 <= lru_127;
      end else begin
        lru_39 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_40 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h28 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_40 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_40 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_40 <= lru_127;
      end else begin
        lru_40 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_41 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h29 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_41 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_41 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_41 <= lru_127;
      end else begin
        lru_41 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_42 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h2a == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_42 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_42 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_42 <= lru_127;
      end else begin
        lru_42 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_43 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h2b == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_43 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_43 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_43 <= lru_127;
      end else begin
        lru_43 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_44 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h2c == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_44 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_44 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_44 <= lru_127;
      end else begin
        lru_44 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_45 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h2d == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_45 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_45 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_45 <= lru_127;
      end else begin
        lru_45 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_46 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h2e == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_46 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_46 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_46 <= lru_127;
      end else begin
        lru_46 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_47 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h2f == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_47 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_47 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_47 <= lru_127;
      end else begin
        lru_47 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_48 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h30 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_48 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_48 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_48 <= lru_127;
      end else begin
        lru_48 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_49 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h31 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_49 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_49 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_49 <= lru_127;
      end else begin
        lru_49 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_50 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h32 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_50 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_50 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_50 <= lru_127;
      end else begin
        lru_50 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_51 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h33 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_51 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_51 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_51 <= lru_127;
      end else begin
        lru_51 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_52 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h34 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_52 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_52 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_52 <= lru_127;
      end else begin
        lru_52 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_53 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h35 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_53 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_53 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_53 <= lru_127;
      end else begin
        lru_53 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_54 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h36 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_54 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_54 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_54 <= lru_127;
      end else begin
        lru_54 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_55 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h37 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_55 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_55 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_55 <= lru_127;
      end else begin
        lru_55 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_56 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h38 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_56 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_56 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_56 <= lru_127;
      end else begin
        lru_56 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_57 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h39 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_57 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_57 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_57 <= lru_127;
      end else begin
        lru_57 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_58 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h3a == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_58 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_58 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_58 <= lru_127;
      end else begin
        lru_58 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_59 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h3b == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_59 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_59 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_59 <= lru_127;
      end else begin
        lru_59 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_60 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h3c == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_60 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_60 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_60 <= lru_127;
      end else begin
        lru_60 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_61 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h3d == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_61 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_61 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_61 <= lru_127;
      end else begin
        lru_61 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_62 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h3e == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_62 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_62 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_62 <= lru_127;
      end else begin
        lru_62 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_63 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h3f == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_63 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_63 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_63 <= lru_127;
      end else begin
        lru_63 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_64 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h40 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_64 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_64 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_64 <= lru_127;
      end else begin
        lru_64 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_65 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h41 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_65 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_65 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_65 <= lru_127;
      end else begin
        lru_65 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_66 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h42 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_66 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_66 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_66 <= lru_127;
      end else begin
        lru_66 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_67 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h43 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_67 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_67 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_67 <= lru_127;
      end else begin
        lru_67 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_68 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h44 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_68 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_68 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_68 <= lru_127;
      end else begin
        lru_68 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_69 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h45 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_69 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_69 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_69 <= lru_127;
      end else begin
        lru_69 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_70 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h46 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_70 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_70 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_70 <= lru_127;
      end else begin
        lru_70 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_71 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h47 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_71 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_71 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_71 <= lru_127;
      end else begin
        lru_71 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_72 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h48 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_72 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_72 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_72 <= lru_127;
      end else begin
        lru_72 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_73 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h49 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_73 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_73 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_73 <= lru_127;
      end else begin
        lru_73 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_74 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h4a == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_74 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_74 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_74 <= lru_127;
      end else begin
        lru_74 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_75 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h4b == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_75 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_75 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_75 <= lru_127;
      end else begin
        lru_75 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_76 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h4c == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_76 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_76 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_76 <= lru_127;
      end else begin
        lru_76 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_77 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h4d == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_77 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_77 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_77 <= lru_127;
      end else begin
        lru_77 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_78 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h4e == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_78 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_78 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_78 <= lru_127;
      end else begin
        lru_78 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_79 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h4f == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_79 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_79 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_79 <= lru_127;
      end else begin
        lru_79 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_80 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h50 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_80 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_80 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_80 <= lru_127;
      end else begin
        lru_80 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_81 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h51 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_81 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_81 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_81 <= lru_127;
      end else begin
        lru_81 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_82 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h52 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_82 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_82 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_82 <= lru_127;
      end else begin
        lru_82 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_83 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h53 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_83 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_83 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_83 <= lru_127;
      end else begin
        lru_83 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_84 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h54 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_84 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_84 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_84 <= lru_127;
      end else begin
        lru_84 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_85 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h55 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_85 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_85 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_85 <= lru_127;
      end else begin
        lru_85 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_86 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h56 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_86 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_86 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_86 <= lru_127;
      end else begin
        lru_86 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_87 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h57 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_87 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_87 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_87 <= lru_127;
      end else begin
        lru_87 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_88 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h58 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_88 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_88 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_88 <= lru_127;
      end else begin
        lru_88 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_89 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h59 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_89 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_89 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_89 <= lru_127;
      end else begin
        lru_89 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_90 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h5a == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_90 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_90 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_90 <= lru_127;
      end else begin
        lru_90 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_91 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h5b == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_91 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_91 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_91 <= lru_127;
      end else begin
        lru_91 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_92 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h5c == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_92 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_92 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_92 <= lru_127;
      end else begin
        lru_92 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_93 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h5d == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_93 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_93 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_93 <= lru_127;
      end else begin
        lru_93 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_94 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h5e == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_94 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_94 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_94 <= lru_127;
      end else begin
        lru_94 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_95 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h5f == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_95 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_95 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_95 <= lru_127;
      end else begin
        lru_95 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_96 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h60 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_96 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_96 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_96 <= lru_127;
      end else begin
        lru_96 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_97 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h61 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_97 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_97 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_97 <= lru_127;
      end else begin
        lru_97 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_98 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h62 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_98 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_98 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_98 <= lru_127;
      end else begin
        lru_98 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_99 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h63 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_99 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_99 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_99 <= lru_127;
      end else begin
        lru_99 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_100 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h64 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_100 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_100 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_100 <= lru_127;
      end else begin
        lru_100 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_101 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h65 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_101 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_101 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_101 <= lru_127;
      end else begin
        lru_101 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_102 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h66 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_102 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_102 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_102 <= lru_127;
      end else begin
        lru_102 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_103 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h67 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_103 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_103 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_103 <= lru_127;
      end else begin
        lru_103 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_104 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h68 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_104 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_104 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_104 <= lru_127;
      end else begin
        lru_104 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_105 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h69 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_105 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_105 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_105 <= lru_127;
      end else begin
        lru_105 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_106 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h6a == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_106 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_106 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_106 <= lru_127;
      end else begin
        lru_106 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_107 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h6b == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_107 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_107 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_107 <= lru_127;
      end else begin
        lru_107 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_108 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h6c == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_108 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_108 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_108 <= lru_127;
      end else begin
        lru_108 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_109 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h6d == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_109 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_109 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_109 <= lru_127;
      end else begin
        lru_109 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_110 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h6e == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_110 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_110 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_110 <= lru_127;
      end else begin
        lru_110 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_111 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h6f == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_111 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_111 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_111 <= lru_127;
      end else begin
        lru_111 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_112 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h70 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_112 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_112 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_112 <= lru_127;
      end else begin
        lru_112 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_113 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h71 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_113 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_113 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_113 <= lru_127;
      end else begin
        lru_113 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_114 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h72 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_114 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_114 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_114 <= lru_127;
      end else begin
        lru_114 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_115 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h73 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_115 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_115 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_115 <= lru_127;
      end else begin
        lru_115 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_116 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h74 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_116 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_116 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_116 <= lru_127;
      end else begin
        lru_116 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_117 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h75 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_117 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_117 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_117 <= lru_127;
      end else begin
        lru_117 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_118 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h76 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_118 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_118 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_118 <= lru_127;
      end else begin
        lru_118 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_119 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h77 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_119 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_119 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_119 <= lru_127;
      end else begin
        lru_119 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_120 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h78 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_120 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_120 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_120 <= lru_127;
      end else begin
        lru_120 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_121 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h79 == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_121 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_121 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_121 <= lru_127;
      end else begin
        lru_121 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_122 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h7a == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_122 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_122 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_122 <= lru_127;
      end else begin
        lru_122 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_123 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h7b == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_123 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_123 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_123 <= lru_127;
      end else begin
        lru_123 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_124 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h7c == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_124 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_124 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_124 <= lru_127;
      end else begin
        lru_124 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_125 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h7d == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_125 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_125 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_125 <= lru_127;
      end else begin
        lru_125 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_126 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h7e == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_126 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_126 <= ~_GEN_130;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_126 <= lru_127;
      end else begin
        lru_126 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 174:37]
      lru_127 <= 1'h0; // @[inst_cache.scala 174:43 176:{12,12} 177:12]
    end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin // @[inst_cache.scala 74:22]
      if (_stage2_stall_T) begin
        lru_127 <= _lru_T_5;
      end else if (_stage1_finished_T_1) begin
        lru_127 <= ~_GEN_130;
      end else if (!(7'h7f == stage1_addr_line_mapping[10:4])) begin
        lru_127 <= _GEN_129;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 244:30]
      work_state <= 4'h1;
    end else if (work_state == 4'h2 & io_port_arready) begin // @[inst_cache.scala 245:12]
      work_state <= 4'h3;
    end else if (_stage1_finished_T_2) begin // @[inst_cache.scala 246:12]
      work_state <= {{1'd0}, _access_work_state_T_7};
    end else if (work_state == 4'h4) begin // @[inst_cache.scala 249:12]
      work_state <= {{1'd0}, _access_work_state_T_22};
    end else if (work_state == 4'h1) begin
      work_state <= {{1'd0}, _access_work_state_T_34};
    end else begin
      work_state <= _access_work_state_T_46;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 264:26]
      write_counter <= 3'h0; // @[inst_cache.scala 264:{106,160}]
    end else if (_access_work_state_T_38 | _stage1_finished_T_2) begin
      if (io_port_rvalid & io_port_rlast) begin
        write_counter <= 3'h0;
      end else if (io_port_rvalid) begin
        write_counter <= _write_counter_T_8;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 258:23]
      wait_data_L <= 40'h0;
    end else if (_stage1_finished_T_2 & io_port_rvalid & _icache_data_way0_0_wen_T_6) begin // @[inst_cache.scala 259:13]
      wait_data_L <= decoder_inst_data;
    end else if (_icache_data_way0_0_wen_T_2 & write_counter == _GEN_1287) begin
      wait_data_L <= decoder_inst_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 110:18 77:28]
      stage1_stall_reg <= 1'h0;
    end else begin
      stage1_stall_reg <= io_sram_req;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      stage1_addr_line_mapping <= 64'h0; // @[inst_cache.scala 118:45]
    end else if (io_sram_req) begin // @[Reg.scala 28:20]
      if (stage1_flush) begin
        stage1_addr_line_mapping <= 64'h0;
      end else begin
        stage1_addr_line_mapping <= io_sram_addr;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 137:38]
      stage1_sram_phy_addr_reg <= 64'h0;
    end else if (stage1_stall_reg) begin
      stage1_sram_phy_addr_reg <= io_p_addr_for_tlb;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      stage1_sram_cache_reg <= 1'h0; // @[inst_cache.scala 120:46]
    end else if (io_sram_req) begin // @[Reg.scala 28:20]
      if (stage1_flush) begin
        stage1_sram_cache_reg <= 1'h0;
      end else begin
        stage1_sram_cache_reg <= io_sram_cache;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      stage1_sram_req_reg <= 1'h0; // @[inst_cache.scala 121:44]
    end else if (_stage1_sram_req_reg_T_1) begin // @[Reg.scala 28:20]
      if (stage1_flush) begin
        stage1_sram_req_reg <= 1'h0;
      end else begin
        stage1_sram_req_reg <= io_inst_ready_to_use;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 140:27]
      stage1_finished <= 1'h0;
    end else if (io_sram_req) begin
      stage1_finished <= 1'h0;
    end else begin
      stage1_finished <= work_state == 4'h7 | work_state == 4'h3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 184:33]
      stage2_sram_addr_reg <= 64'h0;
    end else if (io_stage2_flush) begin // @[inst_cache.scala 184:54]
      stage2_sram_addr_reg <= 64'h0;
    end else if (stage2_stall) begin
      stage2_sram_addr_reg <= stage1_addr_line_mapping;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 190:31]
      stage2_sram_req_reg <= 1'h0;
    end else if (io_stage2_flush) begin // @[inst_cache.scala 190:52]
      stage2_sram_req_reg <= 1'h0;
    end else if (stage2_stall) begin
      stage2_sram_req_reg <= stage1_sram_req_reg;
    end else begin
      stage2_sram_req_reg <= io_sram_write_en == 2'h0 & stage2_sram_req_reg;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 194:27]
      stage2_hit0_reg <= 1'h0;
    end else if (io_stage2_flush) begin // @[inst_cache.scala 194:48]
      stage2_hit0_reg <= 1'h0;
    end else if (stage2_stall) begin
      stage2_hit0_reg <= _hit_T_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 212:31]
      stage2_write_en_reg <= 2'h0;
    end else if (io_stage1_valid_flush) begin // @[inst_cache.scala 212:61]
      stage2_write_en_reg <= 2'h0;
    end else if (stage2_stall) begin
      stage2_write_en_reg <= 2'h1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 145:129]
      has_stage2_stall <= 1'h0;
    end else begin
      has_stage2_stall <= (access_work_state == 4'h1 | access_work_state == 4'h4) & _stage2_stall_T_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[inst_cache.scala 232:28]
      sram_rdata_L_Reg <= 40'h0; // @[inst_cache.scala 221:25 229:{35,84}]
    end else if (has_stage2_stall) begin
      if (_access_work_state_T_8) begin
        sram_rdata_L_Reg <= wait_data_L;
      end else if (_access_work_state_T_23) begin
        if (stage2_hit0_reg) begin
          sram_rdata_L_Reg <= _GEN_516;
        end else begin
          sram_rdata_L_Reg <= _GEN_518;
        end
      end else begin
        sram_rdata_L_Reg <= 40'h0;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  lru_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  lru_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  lru_2 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  lru_3 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  lru_4 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lru_5 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  lru_6 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  lru_7 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  lru_8 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  lru_9 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  lru_10 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  lru_11 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  lru_12 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  lru_13 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  lru_14 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  lru_15 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  lru_16 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  lru_17 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  lru_18 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  lru_19 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  lru_20 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  lru_21 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  lru_22 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  lru_23 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  lru_24 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  lru_25 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  lru_26 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  lru_27 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  lru_28 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  lru_29 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  lru_30 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  lru_31 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  lru_32 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  lru_33 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  lru_34 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  lru_35 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  lru_36 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  lru_37 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  lru_38 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  lru_39 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  lru_40 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  lru_41 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  lru_42 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  lru_43 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  lru_44 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  lru_45 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  lru_46 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  lru_47 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  lru_48 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  lru_49 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  lru_50 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  lru_51 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  lru_52 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  lru_53 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  lru_54 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  lru_55 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  lru_56 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  lru_57 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  lru_58 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  lru_59 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  lru_60 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  lru_61 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  lru_62 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  lru_63 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  lru_64 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  lru_65 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  lru_66 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  lru_67 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  lru_68 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  lru_69 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  lru_70 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  lru_71 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  lru_72 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  lru_73 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  lru_74 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  lru_75 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  lru_76 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  lru_77 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  lru_78 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  lru_79 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  lru_80 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  lru_81 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  lru_82 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  lru_83 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  lru_84 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  lru_85 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  lru_86 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  lru_87 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  lru_88 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  lru_89 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  lru_90 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  lru_91 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  lru_92 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  lru_93 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  lru_94 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  lru_95 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  lru_96 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  lru_97 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  lru_98 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  lru_99 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  lru_100 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  lru_101 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  lru_102 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  lru_103 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  lru_104 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  lru_105 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  lru_106 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  lru_107 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  lru_108 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  lru_109 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  lru_110 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  lru_111 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  lru_112 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  lru_113 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  lru_114 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  lru_115 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  lru_116 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  lru_117 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  lru_118 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  lru_119 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  lru_120 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  lru_121 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  lru_122 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  lru_123 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  lru_124 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  lru_125 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  lru_126 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  lru_127 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  work_state = _RAND_128[3:0];
  _RAND_129 = {1{`RANDOM}};
  write_counter = _RAND_129[2:0];
  _RAND_130 = {2{`RANDOM}};
  wait_data_L = _RAND_130[39:0];
  _RAND_131 = {1{`RANDOM}};
  stage1_stall_reg = _RAND_131[0:0];
  _RAND_132 = {2{`RANDOM}};
  stage1_addr_line_mapping = _RAND_132[63:0];
  _RAND_133 = {2{`RANDOM}};
  stage1_sram_phy_addr_reg = _RAND_133[63:0];
  _RAND_134 = {1{`RANDOM}};
  stage1_sram_cache_reg = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  stage1_sram_req_reg = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  stage1_finished = _RAND_136[0:0];
  _RAND_137 = {2{`RANDOM}};
  stage2_sram_addr_reg = _RAND_137[63:0];
  _RAND_138 = {1{`RANDOM}};
  stage2_sram_req_reg = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  stage2_hit0_reg = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  stage2_write_en_reg = _RAND_140[1:0];
  _RAND_141 = {1{`RANDOM}};
  has_stage2_stall = _RAND_141[0:0];
  _RAND_142 = {2{`RANDOM}};
  sram_rdata_L_Reg = _RAND_142[39:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    lru_0 = 1'h0;
  end
  if (reset) begin
    lru_1 = 1'h0;
  end
  if (reset) begin
    lru_2 = 1'h0;
  end
  if (reset) begin
    lru_3 = 1'h0;
  end
  if (reset) begin
    lru_4 = 1'h0;
  end
  if (reset) begin
    lru_5 = 1'h0;
  end
  if (reset) begin
    lru_6 = 1'h0;
  end
  if (reset) begin
    lru_7 = 1'h0;
  end
  if (reset) begin
    lru_8 = 1'h0;
  end
  if (reset) begin
    lru_9 = 1'h0;
  end
  if (reset) begin
    lru_10 = 1'h0;
  end
  if (reset) begin
    lru_11 = 1'h0;
  end
  if (reset) begin
    lru_12 = 1'h0;
  end
  if (reset) begin
    lru_13 = 1'h0;
  end
  if (reset) begin
    lru_14 = 1'h0;
  end
  if (reset) begin
    lru_15 = 1'h0;
  end
  if (reset) begin
    lru_16 = 1'h0;
  end
  if (reset) begin
    lru_17 = 1'h0;
  end
  if (reset) begin
    lru_18 = 1'h0;
  end
  if (reset) begin
    lru_19 = 1'h0;
  end
  if (reset) begin
    lru_20 = 1'h0;
  end
  if (reset) begin
    lru_21 = 1'h0;
  end
  if (reset) begin
    lru_22 = 1'h0;
  end
  if (reset) begin
    lru_23 = 1'h0;
  end
  if (reset) begin
    lru_24 = 1'h0;
  end
  if (reset) begin
    lru_25 = 1'h0;
  end
  if (reset) begin
    lru_26 = 1'h0;
  end
  if (reset) begin
    lru_27 = 1'h0;
  end
  if (reset) begin
    lru_28 = 1'h0;
  end
  if (reset) begin
    lru_29 = 1'h0;
  end
  if (reset) begin
    lru_30 = 1'h0;
  end
  if (reset) begin
    lru_31 = 1'h0;
  end
  if (reset) begin
    lru_32 = 1'h0;
  end
  if (reset) begin
    lru_33 = 1'h0;
  end
  if (reset) begin
    lru_34 = 1'h0;
  end
  if (reset) begin
    lru_35 = 1'h0;
  end
  if (reset) begin
    lru_36 = 1'h0;
  end
  if (reset) begin
    lru_37 = 1'h0;
  end
  if (reset) begin
    lru_38 = 1'h0;
  end
  if (reset) begin
    lru_39 = 1'h0;
  end
  if (reset) begin
    lru_40 = 1'h0;
  end
  if (reset) begin
    lru_41 = 1'h0;
  end
  if (reset) begin
    lru_42 = 1'h0;
  end
  if (reset) begin
    lru_43 = 1'h0;
  end
  if (reset) begin
    lru_44 = 1'h0;
  end
  if (reset) begin
    lru_45 = 1'h0;
  end
  if (reset) begin
    lru_46 = 1'h0;
  end
  if (reset) begin
    lru_47 = 1'h0;
  end
  if (reset) begin
    lru_48 = 1'h0;
  end
  if (reset) begin
    lru_49 = 1'h0;
  end
  if (reset) begin
    lru_50 = 1'h0;
  end
  if (reset) begin
    lru_51 = 1'h0;
  end
  if (reset) begin
    lru_52 = 1'h0;
  end
  if (reset) begin
    lru_53 = 1'h0;
  end
  if (reset) begin
    lru_54 = 1'h0;
  end
  if (reset) begin
    lru_55 = 1'h0;
  end
  if (reset) begin
    lru_56 = 1'h0;
  end
  if (reset) begin
    lru_57 = 1'h0;
  end
  if (reset) begin
    lru_58 = 1'h0;
  end
  if (reset) begin
    lru_59 = 1'h0;
  end
  if (reset) begin
    lru_60 = 1'h0;
  end
  if (reset) begin
    lru_61 = 1'h0;
  end
  if (reset) begin
    lru_62 = 1'h0;
  end
  if (reset) begin
    lru_63 = 1'h0;
  end
  if (reset) begin
    lru_64 = 1'h0;
  end
  if (reset) begin
    lru_65 = 1'h0;
  end
  if (reset) begin
    lru_66 = 1'h0;
  end
  if (reset) begin
    lru_67 = 1'h0;
  end
  if (reset) begin
    lru_68 = 1'h0;
  end
  if (reset) begin
    lru_69 = 1'h0;
  end
  if (reset) begin
    lru_70 = 1'h0;
  end
  if (reset) begin
    lru_71 = 1'h0;
  end
  if (reset) begin
    lru_72 = 1'h0;
  end
  if (reset) begin
    lru_73 = 1'h0;
  end
  if (reset) begin
    lru_74 = 1'h0;
  end
  if (reset) begin
    lru_75 = 1'h0;
  end
  if (reset) begin
    lru_76 = 1'h0;
  end
  if (reset) begin
    lru_77 = 1'h0;
  end
  if (reset) begin
    lru_78 = 1'h0;
  end
  if (reset) begin
    lru_79 = 1'h0;
  end
  if (reset) begin
    lru_80 = 1'h0;
  end
  if (reset) begin
    lru_81 = 1'h0;
  end
  if (reset) begin
    lru_82 = 1'h0;
  end
  if (reset) begin
    lru_83 = 1'h0;
  end
  if (reset) begin
    lru_84 = 1'h0;
  end
  if (reset) begin
    lru_85 = 1'h0;
  end
  if (reset) begin
    lru_86 = 1'h0;
  end
  if (reset) begin
    lru_87 = 1'h0;
  end
  if (reset) begin
    lru_88 = 1'h0;
  end
  if (reset) begin
    lru_89 = 1'h0;
  end
  if (reset) begin
    lru_90 = 1'h0;
  end
  if (reset) begin
    lru_91 = 1'h0;
  end
  if (reset) begin
    lru_92 = 1'h0;
  end
  if (reset) begin
    lru_93 = 1'h0;
  end
  if (reset) begin
    lru_94 = 1'h0;
  end
  if (reset) begin
    lru_95 = 1'h0;
  end
  if (reset) begin
    lru_96 = 1'h0;
  end
  if (reset) begin
    lru_97 = 1'h0;
  end
  if (reset) begin
    lru_98 = 1'h0;
  end
  if (reset) begin
    lru_99 = 1'h0;
  end
  if (reset) begin
    lru_100 = 1'h0;
  end
  if (reset) begin
    lru_101 = 1'h0;
  end
  if (reset) begin
    lru_102 = 1'h0;
  end
  if (reset) begin
    lru_103 = 1'h0;
  end
  if (reset) begin
    lru_104 = 1'h0;
  end
  if (reset) begin
    lru_105 = 1'h0;
  end
  if (reset) begin
    lru_106 = 1'h0;
  end
  if (reset) begin
    lru_107 = 1'h0;
  end
  if (reset) begin
    lru_108 = 1'h0;
  end
  if (reset) begin
    lru_109 = 1'h0;
  end
  if (reset) begin
    lru_110 = 1'h0;
  end
  if (reset) begin
    lru_111 = 1'h0;
  end
  if (reset) begin
    lru_112 = 1'h0;
  end
  if (reset) begin
    lru_113 = 1'h0;
  end
  if (reset) begin
    lru_114 = 1'h0;
  end
  if (reset) begin
    lru_115 = 1'h0;
  end
  if (reset) begin
    lru_116 = 1'h0;
  end
  if (reset) begin
    lru_117 = 1'h0;
  end
  if (reset) begin
    lru_118 = 1'h0;
  end
  if (reset) begin
    lru_119 = 1'h0;
  end
  if (reset) begin
    lru_120 = 1'h0;
  end
  if (reset) begin
    lru_121 = 1'h0;
  end
  if (reset) begin
    lru_122 = 1'h0;
  end
  if (reset) begin
    lru_123 = 1'h0;
  end
  if (reset) begin
    lru_124 = 1'h0;
  end
  if (reset) begin
    lru_125 = 1'h0;
  end
  if (reset) begin
    lru_126 = 1'h0;
  end
  if (reset) begin
    lru_127 = 1'h0;
  end
  if (reset) begin
    work_state = 4'h1;
  end
  if (reset) begin
    write_counter = 3'h0;
  end
  if (reset) begin
    wait_data_L = 40'h0;
  end
  if (reset) begin
    stage1_stall_reg = 1'h0;
  end
  if (reset) begin
    stage1_addr_line_mapping = 64'h0;
  end
  if (reset) begin
    stage1_sram_phy_addr_reg = 64'h0;
  end
  if (reset) begin
    stage1_sram_cache_reg = 1'h0;
  end
  if (reset) begin
    stage1_sram_req_reg = 1'h0;
  end
  if (reset) begin
    stage1_finished = 1'h0;
  end
  if (reset) begin
    stage2_sram_addr_reg = 64'h0;
  end
  if (reset) begin
    stage2_sram_req_reg = 1'h0;
  end
  if (reset) begin
    stage2_hit0_reg = 1'h0;
  end
  if (reset) begin
    stage2_write_en_reg = 2'h0;
  end
  if (reset) begin
    has_stage2_stall = 1'h0;
  end
  if (reset) begin
    sram_rdata_L_Reg = 40'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module dcache_tag(
  input         clock,
  input         reset,
  input         io_wen,
  input  [53:0] io_wdata,
  input  [63:0] io_raddr,
  input  [63:0] io_waddr,
  output        io_hit,
  output        io_valid,
  output [52:0] io_tag,
  output        io_w_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_43;
  reg [63:0] _RAND_44;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_46;
  reg [63:0] _RAND_47;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_55;
  reg [63:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [63:0] _RAND_62;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_64;
  reg [63:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_67;
  reg [63:0] _RAND_68;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [63:0] _RAND_74;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_76;
  reg [63:0] _RAND_77;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [63:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_82;
  reg [63:0] _RAND_83;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_94;
  reg [63:0] _RAND_95;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_97;
  reg [63:0] _RAND_98;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_103;
  reg [63:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_106;
  reg [63:0] _RAND_107;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_109;
  reg [63:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_112;
  reg [63:0] _RAND_113;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [63:0] _RAND_116;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [63:0] _RAND_119;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [63:0] _RAND_122;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_124;
  reg [63:0] _RAND_125;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_127;
`endif // RANDOMIZE_REG_INIT
  reg [53:0] tag_regs0_0; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_1; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_2; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_3; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_4; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_5; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_6; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_7; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_8; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_9; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_10; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_11; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_12; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_13; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_14; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_15; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_16; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_17; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_18; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_19; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_20; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_21; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_22; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_23; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_24; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_25; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_26; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_27; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_28; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_29; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_30; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_31; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_32; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_33; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_34; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_35; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_36; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_37; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_38; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_39; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_40; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_41; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_42; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_43; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_44; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_45; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_46; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_47; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_48; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_49; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_50; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_51; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_52; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_53; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_54; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_55; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_56; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_57; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_58; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_59; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_60; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_61; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_62; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs0_63; // @[dcache_tag.scala 23:28]
  reg [53:0] tag_regs1_0; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_1; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_2; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_3; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_4; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_5; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_6; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_7; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_8; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_9; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_10; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_11; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_12; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_13; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_14; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_15; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_16; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_17; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_18; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_19; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_20; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_21; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_22; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_23; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_24; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_25; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_26; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_27; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_28; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_29; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_30; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_31; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_32; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_33; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_34; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_35; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_36; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_37; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_38; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_39; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_40; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_41; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_42; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_43; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_44; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_45; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_46; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_47; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_48; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_49; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_50; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_51; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_52; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_53; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_54; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_55; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_56; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_57; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_58; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_59; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_60; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_61; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_62; // @[dcache_tag.scala 24:28]
  reg [53:0] tag_regs1_63; // @[dcache_tag.scala 24:28]
  wire [53:0] _GEN_1 = 6'h1 == io_waddr[10:5] ? tag_regs0_1 : tag_regs0_0; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_2 = 6'h2 == io_waddr[10:5] ? tag_regs0_2 : _GEN_1; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_3 = 6'h3 == io_waddr[10:5] ? tag_regs0_3 : _GEN_2; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_4 = 6'h4 == io_waddr[10:5] ? tag_regs0_4 : _GEN_3; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_5 = 6'h5 == io_waddr[10:5] ? tag_regs0_5 : _GEN_4; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_6 = 6'h6 == io_waddr[10:5] ? tag_regs0_6 : _GEN_5; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_7 = 6'h7 == io_waddr[10:5] ? tag_regs0_7 : _GEN_6; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_8 = 6'h8 == io_waddr[10:5] ? tag_regs0_8 : _GEN_7; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_9 = 6'h9 == io_waddr[10:5] ? tag_regs0_9 : _GEN_8; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_10 = 6'ha == io_waddr[10:5] ? tag_regs0_10 : _GEN_9; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_11 = 6'hb == io_waddr[10:5] ? tag_regs0_11 : _GEN_10; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_12 = 6'hc == io_waddr[10:5] ? tag_regs0_12 : _GEN_11; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_13 = 6'hd == io_waddr[10:5] ? tag_regs0_13 : _GEN_12; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_14 = 6'he == io_waddr[10:5] ? tag_regs0_14 : _GEN_13; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_15 = 6'hf == io_waddr[10:5] ? tag_regs0_15 : _GEN_14; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_16 = 6'h10 == io_waddr[10:5] ? tag_regs0_16 : _GEN_15; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_17 = 6'h11 == io_waddr[10:5] ? tag_regs0_17 : _GEN_16; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_18 = 6'h12 == io_waddr[10:5] ? tag_regs0_18 : _GEN_17; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_19 = 6'h13 == io_waddr[10:5] ? tag_regs0_19 : _GEN_18; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_20 = 6'h14 == io_waddr[10:5] ? tag_regs0_20 : _GEN_19; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_21 = 6'h15 == io_waddr[10:5] ? tag_regs0_21 : _GEN_20; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_22 = 6'h16 == io_waddr[10:5] ? tag_regs0_22 : _GEN_21; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_23 = 6'h17 == io_waddr[10:5] ? tag_regs0_23 : _GEN_22; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_24 = 6'h18 == io_waddr[10:5] ? tag_regs0_24 : _GEN_23; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_25 = 6'h19 == io_waddr[10:5] ? tag_regs0_25 : _GEN_24; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_26 = 6'h1a == io_waddr[10:5] ? tag_regs0_26 : _GEN_25; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_27 = 6'h1b == io_waddr[10:5] ? tag_regs0_27 : _GEN_26; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_28 = 6'h1c == io_waddr[10:5] ? tag_regs0_28 : _GEN_27; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_29 = 6'h1d == io_waddr[10:5] ? tag_regs0_29 : _GEN_28; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_30 = 6'h1e == io_waddr[10:5] ? tag_regs0_30 : _GEN_29; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_31 = 6'h1f == io_waddr[10:5] ? tag_regs0_31 : _GEN_30; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_32 = 6'h20 == io_waddr[10:5] ? tag_regs0_32 : _GEN_31; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_33 = 6'h21 == io_waddr[10:5] ? tag_regs0_33 : _GEN_32; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_34 = 6'h22 == io_waddr[10:5] ? tag_regs0_34 : _GEN_33; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_35 = 6'h23 == io_waddr[10:5] ? tag_regs0_35 : _GEN_34; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_36 = 6'h24 == io_waddr[10:5] ? tag_regs0_36 : _GEN_35; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_37 = 6'h25 == io_waddr[10:5] ? tag_regs0_37 : _GEN_36; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_38 = 6'h26 == io_waddr[10:5] ? tag_regs0_38 : _GEN_37; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_39 = 6'h27 == io_waddr[10:5] ? tag_regs0_39 : _GEN_38; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_40 = 6'h28 == io_waddr[10:5] ? tag_regs0_40 : _GEN_39; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_41 = 6'h29 == io_waddr[10:5] ? tag_regs0_41 : _GEN_40; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_42 = 6'h2a == io_waddr[10:5] ? tag_regs0_42 : _GEN_41; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_43 = 6'h2b == io_waddr[10:5] ? tag_regs0_43 : _GEN_42; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_44 = 6'h2c == io_waddr[10:5] ? tag_regs0_44 : _GEN_43; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_45 = 6'h2d == io_waddr[10:5] ? tag_regs0_45 : _GEN_44; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_46 = 6'h2e == io_waddr[10:5] ? tag_regs0_46 : _GEN_45; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_47 = 6'h2f == io_waddr[10:5] ? tag_regs0_47 : _GEN_46; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_48 = 6'h30 == io_waddr[10:5] ? tag_regs0_48 : _GEN_47; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_49 = 6'h31 == io_waddr[10:5] ? tag_regs0_49 : _GEN_48; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_50 = 6'h32 == io_waddr[10:5] ? tag_regs0_50 : _GEN_49; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_51 = 6'h33 == io_waddr[10:5] ? tag_regs0_51 : _GEN_50; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_52 = 6'h34 == io_waddr[10:5] ? tag_regs0_52 : _GEN_51; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_53 = 6'h35 == io_waddr[10:5] ? tag_regs0_53 : _GEN_52; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_54 = 6'h36 == io_waddr[10:5] ? tag_regs0_54 : _GEN_53; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_55 = 6'h37 == io_waddr[10:5] ? tag_regs0_55 : _GEN_54; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_56 = 6'h38 == io_waddr[10:5] ? tag_regs0_56 : _GEN_55; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_57 = 6'h39 == io_waddr[10:5] ? tag_regs0_57 : _GEN_56; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_58 = 6'h3a == io_waddr[10:5] ? tag_regs0_58 : _GEN_57; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_59 = 6'h3b == io_waddr[10:5] ? tag_regs0_59 : _GEN_58; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_60 = 6'h3c == io_waddr[10:5] ? tag_regs0_60 : _GEN_59; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_61 = 6'h3d == io_waddr[10:5] ? tag_regs0_61 : _GEN_60; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_62 = 6'h3e == io_waddr[10:5] ? tag_regs0_62 : _GEN_61; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_63 = 6'h3f == io_waddr[10:5] ? tag_regs0_63 : _GEN_62; // @[dcache_tag.scala 27:{37,37}]
  wire [53:0] _GEN_129 = 6'h1 == io_waddr[10:5] ? tag_regs1_1 : tag_regs1_0; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_130 = 6'h2 == io_waddr[10:5] ? tag_regs1_2 : _GEN_129; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_131 = 6'h3 == io_waddr[10:5] ? tag_regs1_3 : _GEN_130; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_132 = 6'h4 == io_waddr[10:5] ? tag_regs1_4 : _GEN_131; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_133 = 6'h5 == io_waddr[10:5] ? tag_regs1_5 : _GEN_132; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_134 = 6'h6 == io_waddr[10:5] ? tag_regs1_6 : _GEN_133; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_135 = 6'h7 == io_waddr[10:5] ? tag_regs1_7 : _GEN_134; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_136 = 6'h8 == io_waddr[10:5] ? tag_regs1_8 : _GEN_135; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_137 = 6'h9 == io_waddr[10:5] ? tag_regs1_9 : _GEN_136; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_138 = 6'ha == io_waddr[10:5] ? tag_regs1_10 : _GEN_137; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_139 = 6'hb == io_waddr[10:5] ? tag_regs1_11 : _GEN_138; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_140 = 6'hc == io_waddr[10:5] ? tag_regs1_12 : _GEN_139; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_141 = 6'hd == io_waddr[10:5] ? tag_regs1_13 : _GEN_140; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_142 = 6'he == io_waddr[10:5] ? tag_regs1_14 : _GEN_141; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_143 = 6'hf == io_waddr[10:5] ? tag_regs1_15 : _GEN_142; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_144 = 6'h10 == io_waddr[10:5] ? tag_regs1_16 : _GEN_143; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_145 = 6'h11 == io_waddr[10:5] ? tag_regs1_17 : _GEN_144; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_146 = 6'h12 == io_waddr[10:5] ? tag_regs1_18 : _GEN_145; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_147 = 6'h13 == io_waddr[10:5] ? tag_regs1_19 : _GEN_146; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_148 = 6'h14 == io_waddr[10:5] ? tag_regs1_20 : _GEN_147; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_149 = 6'h15 == io_waddr[10:5] ? tag_regs1_21 : _GEN_148; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_150 = 6'h16 == io_waddr[10:5] ? tag_regs1_22 : _GEN_149; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_151 = 6'h17 == io_waddr[10:5] ? tag_regs1_23 : _GEN_150; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_152 = 6'h18 == io_waddr[10:5] ? tag_regs1_24 : _GEN_151; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_153 = 6'h19 == io_waddr[10:5] ? tag_regs1_25 : _GEN_152; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_154 = 6'h1a == io_waddr[10:5] ? tag_regs1_26 : _GEN_153; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_155 = 6'h1b == io_waddr[10:5] ? tag_regs1_27 : _GEN_154; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_156 = 6'h1c == io_waddr[10:5] ? tag_regs1_28 : _GEN_155; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_157 = 6'h1d == io_waddr[10:5] ? tag_regs1_29 : _GEN_156; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_158 = 6'h1e == io_waddr[10:5] ? tag_regs1_30 : _GEN_157; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_159 = 6'h1f == io_waddr[10:5] ? tag_regs1_31 : _GEN_158; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_160 = 6'h20 == io_waddr[10:5] ? tag_regs1_32 : _GEN_159; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_161 = 6'h21 == io_waddr[10:5] ? tag_regs1_33 : _GEN_160; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_162 = 6'h22 == io_waddr[10:5] ? tag_regs1_34 : _GEN_161; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_163 = 6'h23 == io_waddr[10:5] ? tag_regs1_35 : _GEN_162; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_164 = 6'h24 == io_waddr[10:5] ? tag_regs1_36 : _GEN_163; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_165 = 6'h25 == io_waddr[10:5] ? tag_regs1_37 : _GEN_164; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_166 = 6'h26 == io_waddr[10:5] ? tag_regs1_38 : _GEN_165; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_167 = 6'h27 == io_waddr[10:5] ? tag_regs1_39 : _GEN_166; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_168 = 6'h28 == io_waddr[10:5] ? tag_regs1_40 : _GEN_167; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_169 = 6'h29 == io_waddr[10:5] ? tag_regs1_41 : _GEN_168; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_170 = 6'h2a == io_waddr[10:5] ? tag_regs1_42 : _GEN_169; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_171 = 6'h2b == io_waddr[10:5] ? tag_regs1_43 : _GEN_170; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_172 = 6'h2c == io_waddr[10:5] ? tag_regs1_44 : _GEN_171; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_173 = 6'h2d == io_waddr[10:5] ? tag_regs1_45 : _GEN_172; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_174 = 6'h2e == io_waddr[10:5] ? tag_regs1_46 : _GEN_173; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_175 = 6'h2f == io_waddr[10:5] ? tag_regs1_47 : _GEN_174; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_176 = 6'h30 == io_waddr[10:5] ? tag_regs1_48 : _GEN_175; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_177 = 6'h31 == io_waddr[10:5] ? tag_regs1_49 : _GEN_176; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_178 = 6'h32 == io_waddr[10:5] ? tag_regs1_50 : _GEN_177; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_179 = 6'h33 == io_waddr[10:5] ? tag_regs1_51 : _GEN_178; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_180 = 6'h34 == io_waddr[10:5] ? tag_regs1_52 : _GEN_179; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_181 = 6'h35 == io_waddr[10:5] ? tag_regs1_53 : _GEN_180; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_182 = 6'h36 == io_waddr[10:5] ? tag_regs1_54 : _GEN_181; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_183 = 6'h37 == io_waddr[10:5] ? tag_regs1_55 : _GEN_182; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_184 = 6'h38 == io_waddr[10:5] ? tag_regs1_56 : _GEN_183; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_185 = 6'h39 == io_waddr[10:5] ? tag_regs1_57 : _GEN_184; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_186 = 6'h3a == io_waddr[10:5] ? tag_regs1_58 : _GEN_185; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_187 = 6'h3b == io_waddr[10:5] ? tag_regs1_59 : _GEN_186; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_188 = 6'h3c == io_waddr[10:5] ? tag_regs1_60 : _GEN_187; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_189 = 6'h3d == io_waddr[10:5] ? tag_regs1_61 : _GEN_188; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_190 = 6'h3e == io_waddr[10:5] ? tag_regs1_62 : _GEN_189; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_191 = 6'h3f == io_waddr[10:5] ? tag_regs1_63 : _GEN_190; // @[dcache_tag.scala 28:{37,37}]
  wire [53:0] _GEN_385 = 6'h1 == io_raddr[10:5] ? tag_regs1_1 : tag_regs1_0; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_386 = 6'h2 == io_raddr[10:5] ? tag_regs1_2 : _GEN_385; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_387 = 6'h3 == io_raddr[10:5] ? tag_regs1_3 : _GEN_386; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_388 = 6'h4 == io_raddr[10:5] ? tag_regs1_4 : _GEN_387; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_389 = 6'h5 == io_raddr[10:5] ? tag_regs1_5 : _GEN_388; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_390 = 6'h6 == io_raddr[10:5] ? tag_regs1_6 : _GEN_389; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_391 = 6'h7 == io_raddr[10:5] ? tag_regs1_7 : _GEN_390; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_392 = 6'h8 == io_raddr[10:5] ? tag_regs1_8 : _GEN_391; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_393 = 6'h9 == io_raddr[10:5] ? tag_regs1_9 : _GEN_392; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_394 = 6'ha == io_raddr[10:5] ? tag_regs1_10 : _GEN_393; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_395 = 6'hb == io_raddr[10:5] ? tag_regs1_11 : _GEN_394; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_396 = 6'hc == io_raddr[10:5] ? tag_regs1_12 : _GEN_395; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_397 = 6'hd == io_raddr[10:5] ? tag_regs1_13 : _GEN_396; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_398 = 6'he == io_raddr[10:5] ? tag_regs1_14 : _GEN_397; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_399 = 6'hf == io_raddr[10:5] ? tag_regs1_15 : _GEN_398; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_400 = 6'h10 == io_raddr[10:5] ? tag_regs1_16 : _GEN_399; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_401 = 6'h11 == io_raddr[10:5] ? tag_regs1_17 : _GEN_400; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_402 = 6'h12 == io_raddr[10:5] ? tag_regs1_18 : _GEN_401; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_403 = 6'h13 == io_raddr[10:5] ? tag_regs1_19 : _GEN_402; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_404 = 6'h14 == io_raddr[10:5] ? tag_regs1_20 : _GEN_403; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_405 = 6'h15 == io_raddr[10:5] ? tag_regs1_21 : _GEN_404; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_406 = 6'h16 == io_raddr[10:5] ? tag_regs1_22 : _GEN_405; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_407 = 6'h17 == io_raddr[10:5] ? tag_regs1_23 : _GEN_406; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_408 = 6'h18 == io_raddr[10:5] ? tag_regs1_24 : _GEN_407; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_409 = 6'h19 == io_raddr[10:5] ? tag_regs1_25 : _GEN_408; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_410 = 6'h1a == io_raddr[10:5] ? tag_regs1_26 : _GEN_409; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_411 = 6'h1b == io_raddr[10:5] ? tag_regs1_27 : _GEN_410; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_412 = 6'h1c == io_raddr[10:5] ? tag_regs1_28 : _GEN_411; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_413 = 6'h1d == io_raddr[10:5] ? tag_regs1_29 : _GEN_412; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_414 = 6'h1e == io_raddr[10:5] ? tag_regs1_30 : _GEN_413; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_415 = 6'h1f == io_raddr[10:5] ? tag_regs1_31 : _GEN_414; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_416 = 6'h20 == io_raddr[10:5] ? tag_regs1_32 : _GEN_415; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_417 = 6'h21 == io_raddr[10:5] ? tag_regs1_33 : _GEN_416; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_418 = 6'h22 == io_raddr[10:5] ? tag_regs1_34 : _GEN_417; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_419 = 6'h23 == io_raddr[10:5] ? tag_regs1_35 : _GEN_418; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_420 = 6'h24 == io_raddr[10:5] ? tag_regs1_36 : _GEN_419; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_421 = 6'h25 == io_raddr[10:5] ? tag_regs1_37 : _GEN_420; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_422 = 6'h26 == io_raddr[10:5] ? tag_regs1_38 : _GEN_421; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_423 = 6'h27 == io_raddr[10:5] ? tag_regs1_39 : _GEN_422; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_424 = 6'h28 == io_raddr[10:5] ? tag_regs1_40 : _GEN_423; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_425 = 6'h29 == io_raddr[10:5] ? tag_regs1_41 : _GEN_424; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_426 = 6'h2a == io_raddr[10:5] ? tag_regs1_42 : _GEN_425; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_427 = 6'h2b == io_raddr[10:5] ? tag_regs1_43 : _GEN_426; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_428 = 6'h2c == io_raddr[10:5] ? tag_regs1_44 : _GEN_427; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_429 = 6'h2d == io_raddr[10:5] ? tag_regs1_45 : _GEN_428; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_430 = 6'h2e == io_raddr[10:5] ? tag_regs1_46 : _GEN_429; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_431 = 6'h2f == io_raddr[10:5] ? tag_regs1_47 : _GEN_430; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_432 = 6'h30 == io_raddr[10:5] ? tag_regs1_48 : _GEN_431; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_433 = 6'h31 == io_raddr[10:5] ? tag_regs1_49 : _GEN_432; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_434 = 6'h32 == io_raddr[10:5] ? tag_regs1_50 : _GEN_433; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_435 = 6'h33 == io_raddr[10:5] ? tag_regs1_51 : _GEN_434; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_436 = 6'h34 == io_raddr[10:5] ? tag_regs1_52 : _GEN_435; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_437 = 6'h35 == io_raddr[10:5] ? tag_regs1_53 : _GEN_436; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_438 = 6'h36 == io_raddr[10:5] ? tag_regs1_54 : _GEN_437; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_439 = 6'h37 == io_raddr[10:5] ? tag_regs1_55 : _GEN_438; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_440 = 6'h38 == io_raddr[10:5] ? tag_regs1_56 : _GEN_439; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_441 = 6'h39 == io_raddr[10:5] ? tag_regs1_57 : _GEN_440; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_442 = 6'h3a == io_raddr[10:5] ? tag_regs1_58 : _GEN_441; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_443 = 6'h3b == io_raddr[10:5] ? tag_regs1_59 : _GEN_442; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_444 = 6'h3c == io_raddr[10:5] ? tag_regs1_60 : _GEN_443; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_445 = 6'h3d == io_raddr[10:5] ? tag_regs1_61 : _GEN_444; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_446 = 6'h3e == io_raddr[10:5] ? tag_regs1_62 : _GEN_445; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_447 = 6'h3f == io_raddr[10:5] ? tag_regs1_63 : _GEN_446; // @[dcache_tag.scala 38:{44,44}]
  wire [53:0] _GEN_449 = 6'h1 == io_raddr[10:5] ? tag_regs0_1 : tag_regs0_0; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_450 = 6'h2 == io_raddr[10:5] ? tag_regs0_2 : _GEN_449; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_451 = 6'h3 == io_raddr[10:5] ? tag_regs0_3 : _GEN_450; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_452 = 6'h4 == io_raddr[10:5] ? tag_regs0_4 : _GEN_451; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_453 = 6'h5 == io_raddr[10:5] ? tag_regs0_5 : _GEN_452; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_454 = 6'h6 == io_raddr[10:5] ? tag_regs0_6 : _GEN_453; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_455 = 6'h7 == io_raddr[10:5] ? tag_regs0_7 : _GEN_454; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_456 = 6'h8 == io_raddr[10:5] ? tag_regs0_8 : _GEN_455; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_457 = 6'h9 == io_raddr[10:5] ? tag_regs0_9 : _GEN_456; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_458 = 6'ha == io_raddr[10:5] ? tag_regs0_10 : _GEN_457; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_459 = 6'hb == io_raddr[10:5] ? tag_regs0_11 : _GEN_458; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_460 = 6'hc == io_raddr[10:5] ? tag_regs0_12 : _GEN_459; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_461 = 6'hd == io_raddr[10:5] ? tag_regs0_13 : _GEN_460; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_462 = 6'he == io_raddr[10:5] ? tag_regs0_14 : _GEN_461; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_463 = 6'hf == io_raddr[10:5] ? tag_regs0_15 : _GEN_462; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_464 = 6'h10 == io_raddr[10:5] ? tag_regs0_16 : _GEN_463; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_465 = 6'h11 == io_raddr[10:5] ? tag_regs0_17 : _GEN_464; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_466 = 6'h12 == io_raddr[10:5] ? tag_regs0_18 : _GEN_465; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_467 = 6'h13 == io_raddr[10:5] ? tag_regs0_19 : _GEN_466; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_468 = 6'h14 == io_raddr[10:5] ? tag_regs0_20 : _GEN_467; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_469 = 6'h15 == io_raddr[10:5] ? tag_regs0_21 : _GEN_468; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_470 = 6'h16 == io_raddr[10:5] ? tag_regs0_22 : _GEN_469; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_471 = 6'h17 == io_raddr[10:5] ? tag_regs0_23 : _GEN_470; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_472 = 6'h18 == io_raddr[10:5] ? tag_regs0_24 : _GEN_471; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_473 = 6'h19 == io_raddr[10:5] ? tag_regs0_25 : _GEN_472; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_474 = 6'h1a == io_raddr[10:5] ? tag_regs0_26 : _GEN_473; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_475 = 6'h1b == io_raddr[10:5] ? tag_regs0_27 : _GEN_474; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_476 = 6'h1c == io_raddr[10:5] ? tag_regs0_28 : _GEN_475; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_477 = 6'h1d == io_raddr[10:5] ? tag_regs0_29 : _GEN_476; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_478 = 6'h1e == io_raddr[10:5] ? tag_regs0_30 : _GEN_477; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_479 = 6'h1f == io_raddr[10:5] ? tag_regs0_31 : _GEN_478; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_480 = 6'h20 == io_raddr[10:5] ? tag_regs0_32 : _GEN_479; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_481 = 6'h21 == io_raddr[10:5] ? tag_regs0_33 : _GEN_480; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_482 = 6'h22 == io_raddr[10:5] ? tag_regs0_34 : _GEN_481; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_483 = 6'h23 == io_raddr[10:5] ? tag_regs0_35 : _GEN_482; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_484 = 6'h24 == io_raddr[10:5] ? tag_regs0_36 : _GEN_483; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_485 = 6'h25 == io_raddr[10:5] ? tag_regs0_37 : _GEN_484; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_486 = 6'h26 == io_raddr[10:5] ? tag_regs0_38 : _GEN_485; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_487 = 6'h27 == io_raddr[10:5] ? tag_regs0_39 : _GEN_486; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_488 = 6'h28 == io_raddr[10:5] ? tag_regs0_40 : _GEN_487; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_489 = 6'h29 == io_raddr[10:5] ? tag_regs0_41 : _GEN_488; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_490 = 6'h2a == io_raddr[10:5] ? tag_regs0_42 : _GEN_489; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_491 = 6'h2b == io_raddr[10:5] ? tag_regs0_43 : _GEN_490; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_492 = 6'h2c == io_raddr[10:5] ? tag_regs0_44 : _GEN_491; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_493 = 6'h2d == io_raddr[10:5] ? tag_regs0_45 : _GEN_492; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_494 = 6'h2e == io_raddr[10:5] ? tag_regs0_46 : _GEN_493; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_495 = 6'h2f == io_raddr[10:5] ? tag_regs0_47 : _GEN_494; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_496 = 6'h30 == io_raddr[10:5] ? tag_regs0_48 : _GEN_495; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_497 = 6'h31 == io_raddr[10:5] ? tag_regs0_49 : _GEN_496; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_498 = 6'h32 == io_raddr[10:5] ? tag_regs0_50 : _GEN_497; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_499 = 6'h33 == io_raddr[10:5] ? tag_regs0_51 : _GEN_498; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_500 = 6'h34 == io_raddr[10:5] ? tag_regs0_52 : _GEN_499; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_501 = 6'h35 == io_raddr[10:5] ? tag_regs0_53 : _GEN_500; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_502 = 6'h36 == io_raddr[10:5] ? tag_regs0_54 : _GEN_501; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_503 = 6'h37 == io_raddr[10:5] ? tag_regs0_55 : _GEN_502; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_504 = 6'h38 == io_raddr[10:5] ? tag_regs0_56 : _GEN_503; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_505 = 6'h39 == io_raddr[10:5] ? tag_regs0_57 : _GEN_504; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_506 = 6'h3a == io_raddr[10:5] ? tag_regs0_58 : _GEN_505; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_507 = 6'h3b == io_raddr[10:5] ? tag_regs0_59 : _GEN_506; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_508 = 6'h3c == io_raddr[10:5] ? tag_regs0_60 : _GEN_507; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_509 = 6'h3d == io_raddr[10:5] ? tag_regs0_61 : _GEN_508; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_510 = 6'h3e == io_raddr[10:5] ? tag_regs0_62 : _GEN_509; // @[dcache_tag.scala 38:{68,68}]
  wire [53:0] _GEN_511 = 6'h3f == io_raddr[10:5] ? tag_regs0_63 : _GEN_510; // @[dcache_tag.scala 38:{68,68}]
  assign io_hit = io_raddr[4] & _GEN_447[52:0] == io_raddr[63:11] | ~io_raddr[4] & _GEN_511[52:0] == io_raddr[63:11]; // @[dcache_tag.scala 39:93]
  assign io_valid = io_raddr[4] ? _GEN_447[53] : _GEN_511[53]; // @[dcache_tag.scala 38:20]
  assign io_tag = io_waddr[4] ? _GEN_191[52:0] : _GEN_63[52:0]; // @[dcache_tag.scala 35:18]
  assign io_w_valid = io_waddr[4] ? _GEN_191[53] : _GEN_63[53]; // @[dcache_tag.scala 36:22]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_0 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h0 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_0 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_0 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_0 <= tag_regs0_62;
      end else begin
        tag_regs0_0 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_1 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h1 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_1 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_1 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_1 <= tag_regs0_62;
      end else begin
        tag_regs0_1 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_2 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h2 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_2 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_2 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_2 <= tag_regs0_62;
      end else begin
        tag_regs0_2 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_3 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h3 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_3 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_3 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_3 <= tag_regs0_62;
      end else begin
        tag_regs0_3 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_4 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h4 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_4 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_4 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_4 <= tag_regs0_62;
      end else begin
        tag_regs0_4 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_5 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h5 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_5 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_5 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_5 <= tag_regs0_62;
      end else begin
        tag_regs0_5 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_6 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h6 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_6 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_6 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_6 <= tag_regs0_62;
      end else begin
        tag_regs0_6 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_7 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h7 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_7 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_7 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_7 <= tag_regs0_62;
      end else begin
        tag_regs0_7 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_8 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h8 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_8 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_8 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_8 <= tag_regs0_62;
      end else begin
        tag_regs0_8 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_9 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h9 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_9 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_9 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_9 <= tag_regs0_62;
      end else begin
        tag_regs0_9 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_10 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'ha == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_10 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_10 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_10 <= tag_regs0_62;
      end else begin
        tag_regs0_10 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_11 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'hb == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_11 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_11 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_11 <= tag_regs0_62;
      end else begin
        tag_regs0_11 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_12 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'hc == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_12 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_12 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_12 <= tag_regs0_62;
      end else begin
        tag_regs0_12 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_13 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'hd == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_13 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_13 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_13 <= tag_regs0_62;
      end else begin
        tag_regs0_13 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_14 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'he == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_14 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_14 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_14 <= tag_regs0_62;
      end else begin
        tag_regs0_14 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_15 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'hf == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_15 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_15 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_15 <= tag_regs0_62;
      end else begin
        tag_regs0_15 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_16 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h10 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_16 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_16 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_16 <= tag_regs0_62;
      end else begin
        tag_regs0_16 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_17 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h11 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_17 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_17 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_17 <= tag_regs0_62;
      end else begin
        tag_regs0_17 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_18 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h12 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_18 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_18 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_18 <= tag_regs0_62;
      end else begin
        tag_regs0_18 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_19 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h13 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_19 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_19 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_19 <= tag_regs0_62;
      end else begin
        tag_regs0_19 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_20 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h14 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_20 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_20 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_20 <= tag_regs0_62;
      end else begin
        tag_regs0_20 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_21 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h15 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_21 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_21 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_21 <= tag_regs0_62;
      end else begin
        tag_regs0_21 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_22 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h16 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_22 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_22 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_22 <= tag_regs0_62;
      end else begin
        tag_regs0_22 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_23 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h17 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_23 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_23 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_23 <= tag_regs0_62;
      end else begin
        tag_regs0_23 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_24 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h18 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_24 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_24 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_24 <= tag_regs0_62;
      end else begin
        tag_regs0_24 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_25 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h19 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_25 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_25 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_25 <= tag_regs0_62;
      end else begin
        tag_regs0_25 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_26 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h1a == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_26 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_26 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_26 <= tag_regs0_62;
      end else begin
        tag_regs0_26 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_27 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h1b == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_27 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_27 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_27 <= tag_regs0_62;
      end else begin
        tag_regs0_27 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_28 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h1c == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_28 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_28 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_28 <= tag_regs0_62;
      end else begin
        tag_regs0_28 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_29 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h1d == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_29 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_29 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_29 <= tag_regs0_62;
      end else begin
        tag_regs0_29 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_30 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h1e == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_30 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_30 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_30 <= tag_regs0_62;
      end else begin
        tag_regs0_30 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_31 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h1f == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_31 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_31 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_31 <= tag_regs0_62;
      end else begin
        tag_regs0_31 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_32 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h20 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_32 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_32 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_32 <= tag_regs0_62;
      end else begin
        tag_regs0_32 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_33 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h21 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_33 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_33 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_33 <= tag_regs0_62;
      end else begin
        tag_regs0_33 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_34 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h22 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_34 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_34 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_34 <= tag_regs0_62;
      end else begin
        tag_regs0_34 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_35 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h23 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_35 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_35 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_35 <= tag_regs0_62;
      end else begin
        tag_regs0_35 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_36 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h24 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_36 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_36 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_36 <= tag_regs0_62;
      end else begin
        tag_regs0_36 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_37 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h25 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_37 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_37 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_37 <= tag_regs0_62;
      end else begin
        tag_regs0_37 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_38 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h26 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_38 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_38 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_38 <= tag_regs0_62;
      end else begin
        tag_regs0_38 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_39 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h27 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_39 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_39 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_39 <= tag_regs0_62;
      end else begin
        tag_regs0_39 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_40 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h28 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_40 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_40 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_40 <= tag_regs0_62;
      end else begin
        tag_regs0_40 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_41 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h29 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_41 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_41 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_41 <= tag_regs0_62;
      end else begin
        tag_regs0_41 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_42 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h2a == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_42 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_42 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_42 <= tag_regs0_62;
      end else begin
        tag_regs0_42 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_43 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h2b == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_43 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_43 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_43 <= tag_regs0_62;
      end else begin
        tag_regs0_43 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_44 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h2c == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_44 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_44 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_44 <= tag_regs0_62;
      end else begin
        tag_regs0_44 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_45 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h2d == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_45 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_45 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_45 <= tag_regs0_62;
      end else begin
        tag_regs0_45 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_46 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h2e == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_46 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_46 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_46 <= tag_regs0_62;
      end else begin
        tag_regs0_46 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_47 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h2f == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_47 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_47 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_47 <= tag_regs0_62;
      end else begin
        tag_regs0_47 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_48 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h30 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_48 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_48 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_48 <= tag_regs0_62;
      end else begin
        tag_regs0_48 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_49 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h31 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_49 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_49 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_49 <= tag_regs0_62;
      end else begin
        tag_regs0_49 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_50 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h32 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_50 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_50 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_50 <= tag_regs0_62;
      end else begin
        tag_regs0_50 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_51 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h33 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_51 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_51 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_51 <= tag_regs0_62;
      end else begin
        tag_regs0_51 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_52 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h34 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_52 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_52 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_52 <= tag_regs0_62;
      end else begin
        tag_regs0_52 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_53 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h35 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_53 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_53 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_53 <= tag_regs0_62;
      end else begin
        tag_regs0_53 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_54 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h36 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_54 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_54 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_54 <= tag_regs0_62;
      end else begin
        tag_regs0_54 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_55 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h37 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_55 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_55 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_55 <= tag_regs0_62;
      end else begin
        tag_regs0_55 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_56 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h38 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_56 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_56 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_56 <= tag_regs0_62;
      end else begin
        tag_regs0_56 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_57 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h39 == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_57 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_57 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_57 <= tag_regs0_62;
      end else begin
        tag_regs0_57 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_58 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h3a == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_58 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_58 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_58 <= tag_regs0_62;
      end else begin
        tag_regs0_58 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_59 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h3b == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_59 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_59 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_59 <= tag_regs0_62;
      end else begin
        tag_regs0_59 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_60 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h3c == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_60 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_60 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_60 <= tag_regs0_62;
      end else begin
        tag_regs0_60 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_61 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h3d == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_61 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_61 <= tag_regs0_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs0_61 <= tag_regs0_62;
      end else begin
        tag_regs0_61 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_62 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h3e == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_62 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs0_62 <= tag_regs0_63;
      end else if (!(6'h3e == io_waddr[10:5])) begin
        tag_regs0_62 <= _GEN_61;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 27:31]
      tag_regs0_63 <= 54'h0; // @[dcache_tag.scala 27:{37,37,37,37,37}]
    end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 23:28]
      if (io_wen & ~io_waddr[4]) begin
        tag_regs0_63 <= io_wdata;
      end else if (!(6'h3f == io_waddr[10:5])) begin
        if (6'h3e == io_waddr[10:5]) begin
          tag_regs0_63 <= tag_regs0_62;
        end else begin
          tag_regs0_63 <= _GEN_61;
        end
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_0 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h0 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_0 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_0 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_0 <= tag_regs1_62;
      end else begin
        tag_regs1_0 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_1 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h1 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_1 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_1 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_1 <= tag_regs1_62;
      end else begin
        tag_regs1_1 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_2 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h2 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_2 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_2 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_2 <= tag_regs1_62;
      end else begin
        tag_regs1_2 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_3 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h3 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_3 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_3 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_3 <= tag_regs1_62;
      end else begin
        tag_regs1_3 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_4 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h4 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_4 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_4 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_4 <= tag_regs1_62;
      end else begin
        tag_regs1_4 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_5 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h5 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_5 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_5 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_5 <= tag_regs1_62;
      end else begin
        tag_regs1_5 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_6 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h6 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_6 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_6 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_6 <= tag_regs1_62;
      end else begin
        tag_regs1_6 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_7 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h7 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_7 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_7 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_7 <= tag_regs1_62;
      end else begin
        tag_regs1_7 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_8 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h8 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_8 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_8 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_8 <= tag_regs1_62;
      end else begin
        tag_regs1_8 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_9 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h9 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_9 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_9 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_9 <= tag_regs1_62;
      end else begin
        tag_regs1_9 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_10 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'ha == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_10 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_10 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_10 <= tag_regs1_62;
      end else begin
        tag_regs1_10 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_11 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'hb == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_11 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_11 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_11 <= tag_regs1_62;
      end else begin
        tag_regs1_11 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_12 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'hc == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_12 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_12 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_12 <= tag_regs1_62;
      end else begin
        tag_regs1_12 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_13 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'hd == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_13 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_13 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_13 <= tag_regs1_62;
      end else begin
        tag_regs1_13 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_14 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'he == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_14 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_14 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_14 <= tag_regs1_62;
      end else begin
        tag_regs1_14 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_15 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'hf == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_15 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_15 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_15 <= tag_regs1_62;
      end else begin
        tag_regs1_15 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_16 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h10 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_16 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_16 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_16 <= tag_regs1_62;
      end else begin
        tag_regs1_16 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_17 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h11 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_17 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_17 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_17 <= tag_regs1_62;
      end else begin
        tag_regs1_17 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_18 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h12 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_18 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_18 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_18 <= tag_regs1_62;
      end else begin
        tag_regs1_18 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_19 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h13 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_19 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_19 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_19 <= tag_regs1_62;
      end else begin
        tag_regs1_19 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_20 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h14 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_20 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_20 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_20 <= tag_regs1_62;
      end else begin
        tag_regs1_20 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_21 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h15 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_21 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_21 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_21 <= tag_regs1_62;
      end else begin
        tag_regs1_21 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_22 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h16 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_22 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_22 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_22 <= tag_regs1_62;
      end else begin
        tag_regs1_22 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_23 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h17 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_23 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_23 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_23 <= tag_regs1_62;
      end else begin
        tag_regs1_23 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_24 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h18 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_24 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_24 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_24 <= tag_regs1_62;
      end else begin
        tag_regs1_24 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_25 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h19 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_25 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_25 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_25 <= tag_regs1_62;
      end else begin
        tag_regs1_25 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_26 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h1a == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_26 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_26 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_26 <= tag_regs1_62;
      end else begin
        tag_regs1_26 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_27 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h1b == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_27 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_27 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_27 <= tag_regs1_62;
      end else begin
        tag_regs1_27 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_28 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h1c == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_28 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_28 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_28 <= tag_regs1_62;
      end else begin
        tag_regs1_28 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_29 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h1d == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_29 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_29 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_29 <= tag_regs1_62;
      end else begin
        tag_regs1_29 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_30 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h1e == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_30 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_30 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_30 <= tag_regs1_62;
      end else begin
        tag_regs1_30 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_31 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h1f == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_31 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_31 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_31 <= tag_regs1_62;
      end else begin
        tag_regs1_31 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_32 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h20 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_32 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_32 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_32 <= tag_regs1_62;
      end else begin
        tag_regs1_32 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_33 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h21 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_33 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_33 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_33 <= tag_regs1_62;
      end else begin
        tag_regs1_33 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_34 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h22 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_34 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_34 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_34 <= tag_regs1_62;
      end else begin
        tag_regs1_34 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_35 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h23 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_35 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_35 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_35 <= tag_regs1_62;
      end else begin
        tag_regs1_35 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_36 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h24 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_36 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_36 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_36 <= tag_regs1_62;
      end else begin
        tag_regs1_36 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_37 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h25 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_37 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_37 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_37 <= tag_regs1_62;
      end else begin
        tag_regs1_37 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_38 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h26 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_38 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_38 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_38 <= tag_regs1_62;
      end else begin
        tag_regs1_38 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_39 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h27 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_39 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_39 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_39 <= tag_regs1_62;
      end else begin
        tag_regs1_39 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_40 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h28 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_40 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_40 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_40 <= tag_regs1_62;
      end else begin
        tag_regs1_40 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_41 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h29 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_41 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_41 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_41 <= tag_regs1_62;
      end else begin
        tag_regs1_41 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_42 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h2a == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_42 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_42 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_42 <= tag_regs1_62;
      end else begin
        tag_regs1_42 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_43 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h2b == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_43 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_43 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_43 <= tag_regs1_62;
      end else begin
        tag_regs1_43 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_44 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h2c == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_44 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_44 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_44 <= tag_regs1_62;
      end else begin
        tag_regs1_44 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_45 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h2d == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_45 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_45 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_45 <= tag_regs1_62;
      end else begin
        tag_regs1_45 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_46 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h2e == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_46 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_46 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_46 <= tag_regs1_62;
      end else begin
        tag_regs1_46 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_47 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h2f == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_47 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_47 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_47 <= tag_regs1_62;
      end else begin
        tag_regs1_47 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_48 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h30 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_48 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_48 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_48 <= tag_regs1_62;
      end else begin
        tag_regs1_48 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_49 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h31 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_49 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_49 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_49 <= tag_regs1_62;
      end else begin
        tag_regs1_49 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_50 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h32 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_50 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_50 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_50 <= tag_regs1_62;
      end else begin
        tag_regs1_50 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_51 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h33 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_51 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_51 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_51 <= tag_regs1_62;
      end else begin
        tag_regs1_51 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_52 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h34 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_52 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_52 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_52 <= tag_regs1_62;
      end else begin
        tag_regs1_52 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_53 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h35 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_53 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_53 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_53 <= tag_regs1_62;
      end else begin
        tag_regs1_53 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_54 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h36 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_54 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_54 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_54 <= tag_regs1_62;
      end else begin
        tag_regs1_54 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_55 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h37 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_55 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_55 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_55 <= tag_regs1_62;
      end else begin
        tag_regs1_55 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_56 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h38 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_56 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_56 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_56 <= tag_regs1_62;
      end else begin
        tag_regs1_56 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_57 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h39 == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_57 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_57 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_57 <= tag_regs1_62;
      end else begin
        tag_regs1_57 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_58 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h3a == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_58 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_58 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_58 <= tag_regs1_62;
      end else begin
        tag_regs1_58 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_59 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h3b == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_59 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_59 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_59 <= tag_regs1_62;
      end else begin
        tag_regs1_59 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_60 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h3c == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_60 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_60 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_60 <= tag_regs1_62;
      end else begin
        tag_regs1_60 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_61 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h3d == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_61 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_61 <= tag_regs1_63;
      end else if (6'h3e == io_waddr[10:5]) begin
        tag_regs1_61 <= tag_regs1_62;
      end else begin
        tag_regs1_61 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_62 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h3e == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_62 <= io_wdata;
      end else if (6'h3f == io_waddr[10:5]) begin
        tag_regs1_62 <= tag_regs1_63;
      end else if (!(6'h3e == io_waddr[10:5])) begin
        tag_regs1_62 <= _GEN_189;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[dcache_tag.scala 28:31]
      tag_regs1_63 <= 54'h0; // @[dcache_tag.scala 28:{37,37,37,37,37}]
    end else if (6'h3f == io_waddr[10:5]) begin // @[dcache_tag.scala 24:28]
      if (io_wen & io_waddr[4]) begin
        tag_regs1_63 <= io_wdata;
      end else if (!(6'h3f == io_waddr[10:5])) begin
        if (6'h3e == io_waddr[10:5]) begin
          tag_regs1_63 <= tag_regs1_62;
        end else begin
          tag_regs1_63 <= _GEN_189;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  tag_regs0_0 = _RAND_0[53:0];
  _RAND_1 = {2{`RANDOM}};
  tag_regs0_1 = _RAND_1[53:0];
  _RAND_2 = {2{`RANDOM}};
  tag_regs0_2 = _RAND_2[53:0];
  _RAND_3 = {2{`RANDOM}};
  tag_regs0_3 = _RAND_3[53:0];
  _RAND_4 = {2{`RANDOM}};
  tag_regs0_4 = _RAND_4[53:0];
  _RAND_5 = {2{`RANDOM}};
  tag_regs0_5 = _RAND_5[53:0];
  _RAND_6 = {2{`RANDOM}};
  tag_regs0_6 = _RAND_6[53:0];
  _RAND_7 = {2{`RANDOM}};
  tag_regs0_7 = _RAND_7[53:0];
  _RAND_8 = {2{`RANDOM}};
  tag_regs0_8 = _RAND_8[53:0];
  _RAND_9 = {2{`RANDOM}};
  tag_regs0_9 = _RAND_9[53:0];
  _RAND_10 = {2{`RANDOM}};
  tag_regs0_10 = _RAND_10[53:0];
  _RAND_11 = {2{`RANDOM}};
  tag_regs0_11 = _RAND_11[53:0];
  _RAND_12 = {2{`RANDOM}};
  tag_regs0_12 = _RAND_12[53:0];
  _RAND_13 = {2{`RANDOM}};
  tag_regs0_13 = _RAND_13[53:0];
  _RAND_14 = {2{`RANDOM}};
  tag_regs0_14 = _RAND_14[53:0];
  _RAND_15 = {2{`RANDOM}};
  tag_regs0_15 = _RAND_15[53:0];
  _RAND_16 = {2{`RANDOM}};
  tag_regs0_16 = _RAND_16[53:0];
  _RAND_17 = {2{`RANDOM}};
  tag_regs0_17 = _RAND_17[53:0];
  _RAND_18 = {2{`RANDOM}};
  tag_regs0_18 = _RAND_18[53:0];
  _RAND_19 = {2{`RANDOM}};
  tag_regs0_19 = _RAND_19[53:0];
  _RAND_20 = {2{`RANDOM}};
  tag_regs0_20 = _RAND_20[53:0];
  _RAND_21 = {2{`RANDOM}};
  tag_regs0_21 = _RAND_21[53:0];
  _RAND_22 = {2{`RANDOM}};
  tag_regs0_22 = _RAND_22[53:0];
  _RAND_23 = {2{`RANDOM}};
  tag_regs0_23 = _RAND_23[53:0];
  _RAND_24 = {2{`RANDOM}};
  tag_regs0_24 = _RAND_24[53:0];
  _RAND_25 = {2{`RANDOM}};
  tag_regs0_25 = _RAND_25[53:0];
  _RAND_26 = {2{`RANDOM}};
  tag_regs0_26 = _RAND_26[53:0];
  _RAND_27 = {2{`RANDOM}};
  tag_regs0_27 = _RAND_27[53:0];
  _RAND_28 = {2{`RANDOM}};
  tag_regs0_28 = _RAND_28[53:0];
  _RAND_29 = {2{`RANDOM}};
  tag_regs0_29 = _RAND_29[53:0];
  _RAND_30 = {2{`RANDOM}};
  tag_regs0_30 = _RAND_30[53:0];
  _RAND_31 = {2{`RANDOM}};
  tag_regs0_31 = _RAND_31[53:0];
  _RAND_32 = {2{`RANDOM}};
  tag_regs0_32 = _RAND_32[53:0];
  _RAND_33 = {2{`RANDOM}};
  tag_regs0_33 = _RAND_33[53:0];
  _RAND_34 = {2{`RANDOM}};
  tag_regs0_34 = _RAND_34[53:0];
  _RAND_35 = {2{`RANDOM}};
  tag_regs0_35 = _RAND_35[53:0];
  _RAND_36 = {2{`RANDOM}};
  tag_regs0_36 = _RAND_36[53:0];
  _RAND_37 = {2{`RANDOM}};
  tag_regs0_37 = _RAND_37[53:0];
  _RAND_38 = {2{`RANDOM}};
  tag_regs0_38 = _RAND_38[53:0];
  _RAND_39 = {2{`RANDOM}};
  tag_regs0_39 = _RAND_39[53:0];
  _RAND_40 = {2{`RANDOM}};
  tag_regs0_40 = _RAND_40[53:0];
  _RAND_41 = {2{`RANDOM}};
  tag_regs0_41 = _RAND_41[53:0];
  _RAND_42 = {2{`RANDOM}};
  tag_regs0_42 = _RAND_42[53:0];
  _RAND_43 = {2{`RANDOM}};
  tag_regs0_43 = _RAND_43[53:0];
  _RAND_44 = {2{`RANDOM}};
  tag_regs0_44 = _RAND_44[53:0];
  _RAND_45 = {2{`RANDOM}};
  tag_regs0_45 = _RAND_45[53:0];
  _RAND_46 = {2{`RANDOM}};
  tag_regs0_46 = _RAND_46[53:0];
  _RAND_47 = {2{`RANDOM}};
  tag_regs0_47 = _RAND_47[53:0];
  _RAND_48 = {2{`RANDOM}};
  tag_regs0_48 = _RAND_48[53:0];
  _RAND_49 = {2{`RANDOM}};
  tag_regs0_49 = _RAND_49[53:0];
  _RAND_50 = {2{`RANDOM}};
  tag_regs0_50 = _RAND_50[53:0];
  _RAND_51 = {2{`RANDOM}};
  tag_regs0_51 = _RAND_51[53:0];
  _RAND_52 = {2{`RANDOM}};
  tag_regs0_52 = _RAND_52[53:0];
  _RAND_53 = {2{`RANDOM}};
  tag_regs0_53 = _RAND_53[53:0];
  _RAND_54 = {2{`RANDOM}};
  tag_regs0_54 = _RAND_54[53:0];
  _RAND_55 = {2{`RANDOM}};
  tag_regs0_55 = _RAND_55[53:0];
  _RAND_56 = {2{`RANDOM}};
  tag_regs0_56 = _RAND_56[53:0];
  _RAND_57 = {2{`RANDOM}};
  tag_regs0_57 = _RAND_57[53:0];
  _RAND_58 = {2{`RANDOM}};
  tag_regs0_58 = _RAND_58[53:0];
  _RAND_59 = {2{`RANDOM}};
  tag_regs0_59 = _RAND_59[53:0];
  _RAND_60 = {2{`RANDOM}};
  tag_regs0_60 = _RAND_60[53:0];
  _RAND_61 = {2{`RANDOM}};
  tag_regs0_61 = _RAND_61[53:0];
  _RAND_62 = {2{`RANDOM}};
  tag_regs0_62 = _RAND_62[53:0];
  _RAND_63 = {2{`RANDOM}};
  tag_regs0_63 = _RAND_63[53:0];
  _RAND_64 = {2{`RANDOM}};
  tag_regs1_0 = _RAND_64[53:0];
  _RAND_65 = {2{`RANDOM}};
  tag_regs1_1 = _RAND_65[53:0];
  _RAND_66 = {2{`RANDOM}};
  tag_regs1_2 = _RAND_66[53:0];
  _RAND_67 = {2{`RANDOM}};
  tag_regs1_3 = _RAND_67[53:0];
  _RAND_68 = {2{`RANDOM}};
  tag_regs1_4 = _RAND_68[53:0];
  _RAND_69 = {2{`RANDOM}};
  tag_regs1_5 = _RAND_69[53:0];
  _RAND_70 = {2{`RANDOM}};
  tag_regs1_6 = _RAND_70[53:0];
  _RAND_71 = {2{`RANDOM}};
  tag_regs1_7 = _RAND_71[53:0];
  _RAND_72 = {2{`RANDOM}};
  tag_regs1_8 = _RAND_72[53:0];
  _RAND_73 = {2{`RANDOM}};
  tag_regs1_9 = _RAND_73[53:0];
  _RAND_74 = {2{`RANDOM}};
  tag_regs1_10 = _RAND_74[53:0];
  _RAND_75 = {2{`RANDOM}};
  tag_regs1_11 = _RAND_75[53:0];
  _RAND_76 = {2{`RANDOM}};
  tag_regs1_12 = _RAND_76[53:0];
  _RAND_77 = {2{`RANDOM}};
  tag_regs1_13 = _RAND_77[53:0];
  _RAND_78 = {2{`RANDOM}};
  tag_regs1_14 = _RAND_78[53:0];
  _RAND_79 = {2{`RANDOM}};
  tag_regs1_15 = _RAND_79[53:0];
  _RAND_80 = {2{`RANDOM}};
  tag_regs1_16 = _RAND_80[53:0];
  _RAND_81 = {2{`RANDOM}};
  tag_regs1_17 = _RAND_81[53:0];
  _RAND_82 = {2{`RANDOM}};
  tag_regs1_18 = _RAND_82[53:0];
  _RAND_83 = {2{`RANDOM}};
  tag_regs1_19 = _RAND_83[53:0];
  _RAND_84 = {2{`RANDOM}};
  tag_regs1_20 = _RAND_84[53:0];
  _RAND_85 = {2{`RANDOM}};
  tag_regs1_21 = _RAND_85[53:0];
  _RAND_86 = {2{`RANDOM}};
  tag_regs1_22 = _RAND_86[53:0];
  _RAND_87 = {2{`RANDOM}};
  tag_regs1_23 = _RAND_87[53:0];
  _RAND_88 = {2{`RANDOM}};
  tag_regs1_24 = _RAND_88[53:0];
  _RAND_89 = {2{`RANDOM}};
  tag_regs1_25 = _RAND_89[53:0];
  _RAND_90 = {2{`RANDOM}};
  tag_regs1_26 = _RAND_90[53:0];
  _RAND_91 = {2{`RANDOM}};
  tag_regs1_27 = _RAND_91[53:0];
  _RAND_92 = {2{`RANDOM}};
  tag_regs1_28 = _RAND_92[53:0];
  _RAND_93 = {2{`RANDOM}};
  tag_regs1_29 = _RAND_93[53:0];
  _RAND_94 = {2{`RANDOM}};
  tag_regs1_30 = _RAND_94[53:0];
  _RAND_95 = {2{`RANDOM}};
  tag_regs1_31 = _RAND_95[53:0];
  _RAND_96 = {2{`RANDOM}};
  tag_regs1_32 = _RAND_96[53:0];
  _RAND_97 = {2{`RANDOM}};
  tag_regs1_33 = _RAND_97[53:0];
  _RAND_98 = {2{`RANDOM}};
  tag_regs1_34 = _RAND_98[53:0];
  _RAND_99 = {2{`RANDOM}};
  tag_regs1_35 = _RAND_99[53:0];
  _RAND_100 = {2{`RANDOM}};
  tag_regs1_36 = _RAND_100[53:0];
  _RAND_101 = {2{`RANDOM}};
  tag_regs1_37 = _RAND_101[53:0];
  _RAND_102 = {2{`RANDOM}};
  tag_regs1_38 = _RAND_102[53:0];
  _RAND_103 = {2{`RANDOM}};
  tag_regs1_39 = _RAND_103[53:0];
  _RAND_104 = {2{`RANDOM}};
  tag_regs1_40 = _RAND_104[53:0];
  _RAND_105 = {2{`RANDOM}};
  tag_regs1_41 = _RAND_105[53:0];
  _RAND_106 = {2{`RANDOM}};
  tag_regs1_42 = _RAND_106[53:0];
  _RAND_107 = {2{`RANDOM}};
  tag_regs1_43 = _RAND_107[53:0];
  _RAND_108 = {2{`RANDOM}};
  tag_regs1_44 = _RAND_108[53:0];
  _RAND_109 = {2{`RANDOM}};
  tag_regs1_45 = _RAND_109[53:0];
  _RAND_110 = {2{`RANDOM}};
  tag_regs1_46 = _RAND_110[53:0];
  _RAND_111 = {2{`RANDOM}};
  tag_regs1_47 = _RAND_111[53:0];
  _RAND_112 = {2{`RANDOM}};
  tag_regs1_48 = _RAND_112[53:0];
  _RAND_113 = {2{`RANDOM}};
  tag_regs1_49 = _RAND_113[53:0];
  _RAND_114 = {2{`RANDOM}};
  tag_regs1_50 = _RAND_114[53:0];
  _RAND_115 = {2{`RANDOM}};
  tag_regs1_51 = _RAND_115[53:0];
  _RAND_116 = {2{`RANDOM}};
  tag_regs1_52 = _RAND_116[53:0];
  _RAND_117 = {2{`RANDOM}};
  tag_regs1_53 = _RAND_117[53:0];
  _RAND_118 = {2{`RANDOM}};
  tag_regs1_54 = _RAND_118[53:0];
  _RAND_119 = {2{`RANDOM}};
  tag_regs1_55 = _RAND_119[53:0];
  _RAND_120 = {2{`RANDOM}};
  tag_regs1_56 = _RAND_120[53:0];
  _RAND_121 = {2{`RANDOM}};
  tag_regs1_57 = _RAND_121[53:0];
  _RAND_122 = {2{`RANDOM}};
  tag_regs1_58 = _RAND_122[53:0];
  _RAND_123 = {2{`RANDOM}};
  tag_regs1_59 = _RAND_123[53:0];
  _RAND_124 = {2{`RANDOM}};
  tag_regs1_60 = _RAND_124[53:0];
  _RAND_125 = {2{`RANDOM}};
  tag_regs1_61 = _RAND_125[53:0];
  _RAND_126 = {2{`RANDOM}};
  tag_regs1_62 = _RAND_126[53:0];
  _RAND_127 = {2{`RANDOM}};
  tag_regs1_63 = _RAND_127[53:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    tag_regs0_0 = 54'h0;
  end
  if (reset) begin
    tag_regs0_1 = 54'h0;
  end
  if (reset) begin
    tag_regs0_2 = 54'h0;
  end
  if (reset) begin
    tag_regs0_3 = 54'h0;
  end
  if (reset) begin
    tag_regs0_4 = 54'h0;
  end
  if (reset) begin
    tag_regs0_5 = 54'h0;
  end
  if (reset) begin
    tag_regs0_6 = 54'h0;
  end
  if (reset) begin
    tag_regs0_7 = 54'h0;
  end
  if (reset) begin
    tag_regs0_8 = 54'h0;
  end
  if (reset) begin
    tag_regs0_9 = 54'h0;
  end
  if (reset) begin
    tag_regs0_10 = 54'h0;
  end
  if (reset) begin
    tag_regs0_11 = 54'h0;
  end
  if (reset) begin
    tag_regs0_12 = 54'h0;
  end
  if (reset) begin
    tag_regs0_13 = 54'h0;
  end
  if (reset) begin
    tag_regs0_14 = 54'h0;
  end
  if (reset) begin
    tag_regs0_15 = 54'h0;
  end
  if (reset) begin
    tag_regs0_16 = 54'h0;
  end
  if (reset) begin
    tag_regs0_17 = 54'h0;
  end
  if (reset) begin
    tag_regs0_18 = 54'h0;
  end
  if (reset) begin
    tag_regs0_19 = 54'h0;
  end
  if (reset) begin
    tag_regs0_20 = 54'h0;
  end
  if (reset) begin
    tag_regs0_21 = 54'h0;
  end
  if (reset) begin
    tag_regs0_22 = 54'h0;
  end
  if (reset) begin
    tag_regs0_23 = 54'h0;
  end
  if (reset) begin
    tag_regs0_24 = 54'h0;
  end
  if (reset) begin
    tag_regs0_25 = 54'h0;
  end
  if (reset) begin
    tag_regs0_26 = 54'h0;
  end
  if (reset) begin
    tag_regs0_27 = 54'h0;
  end
  if (reset) begin
    tag_regs0_28 = 54'h0;
  end
  if (reset) begin
    tag_regs0_29 = 54'h0;
  end
  if (reset) begin
    tag_regs0_30 = 54'h0;
  end
  if (reset) begin
    tag_regs0_31 = 54'h0;
  end
  if (reset) begin
    tag_regs0_32 = 54'h0;
  end
  if (reset) begin
    tag_regs0_33 = 54'h0;
  end
  if (reset) begin
    tag_regs0_34 = 54'h0;
  end
  if (reset) begin
    tag_regs0_35 = 54'h0;
  end
  if (reset) begin
    tag_regs0_36 = 54'h0;
  end
  if (reset) begin
    tag_regs0_37 = 54'h0;
  end
  if (reset) begin
    tag_regs0_38 = 54'h0;
  end
  if (reset) begin
    tag_regs0_39 = 54'h0;
  end
  if (reset) begin
    tag_regs0_40 = 54'h0;
  end
  if (reset) begin
    tag_regs0_41 = 54'h0;
  end
  if (reset) begin
    tag_regs0_42 = 54'h0;
  end
  if (reset) begin
    tag_regs0_43 = 54'h0;
  end
  if (reset) begin
    tag_regs0_44 = 54'h0;
  end
  if (reset) begin
    tag_regs0_45 = 54'h0;
  end
  if (reset) begin
    tag_regs0_46 = 54'h0;
  end
  if (reset) begin
    tag_regs0_47 = 54'h0;
  end
  if (reset) begin
    tag_regs0_48 = 54'h0;
  end
  if (reset) begin
    tag_regs0_49 = 54'h0;
  end
  if (reset) begin
    tag_regs0_50 = 54'h0;
  end
  if (reset) begin
    tag_regs0_51 = 54'h0;
  end
  if (reset) begin
    tag_regs0_52 = 54'h0;
  end
  if (reset) begin
    tag_regs0_53 = 54'h0;
  end
  if (reset) begin
    tag_regs0_54 = 54'h0;
  end
  if (reset) begin
    tag_regs0_55 = 54'h0;
  end
  if (reset) begin
    tag_regs0_56 = 54'h0;
  end
  if (reset) begin
    tag_regs0_57 = 54'h0;
  end
  if (reset) begin
    tag_regs0_58 = 54'h0;
  end
  if (reset) begin
    tag_regs0_59 = 54'h0;
  end
  if (reset) begin
    tag_regs0_60 = 54'h0;
  end
  if (reset) begin
    tag_regs0_61 = 54'h0;
  end
  if (reset) begin
    tag_regs0_62 = 54'h0;
  end
  if (reset) begin
    tag_regs0_63 = 54'h0;
  end
  if (reset) begin
    tag_regs1_0 = 54'h0;
  end
  if (reset) begin
    tag_regs1_1 = 54'h0;
  end
  if (reset) begin
    tag_regs1_2 = 54'h0;
  end
  if (reset) begin
    tag_regs1_3 = 54'h0;
  end
  if (reset) begin
    tag_regs1_4 = 54'h0;
  end
  if (reset) begin
    tag_regs1_5 = 54'h0;
  end
  if (reset) begin
    tag_regs1_6 = 54'h0;
  end
  if (reset) begin
    tag_regs1_7 = 54'h0;
  end
  if (reset) begin
    tag_regs1_8 = 54'h0;
  end
  if (reset) begin
    tag_regs1_9 = 54'h0;
  end
  if (reset) begin
    tag_regs1_10 = 54'h0;
  end
  if (reset) begin
    tag_regs1_11 = 54'h0;
  end
  if (reset) begin
    tag_regs1_12 = 54'h0;
  end
  if (reset) begin
    tag_regs1_13 = 54'h0;
  end
  if (reset) begin
    tag_regs1_14 = 54'h0;
  end
  if (reset) begin
    tag_regs1_15 = 54'h0;
  end
  if (reset) begin
    tag_regs1_16 = 54'h0;
  end
  if (reset) begin
    tag_regs1_17 = 54'h0;
  end
  if (reset) begin
    tag_regs1_18 = 54'h0;
  end
  if (reset) begin
    tag_regs1_19 = 54'h0;
  end
  if (reset) begin
    tag_regs1_20 = 54'h0;
  end
  if (reset) begin
    tag_regs1_21 = 54'h0;
  end
  if (reset) begin
    tag_regs1_22 = 54'h0;
  end
  if (reset) begin
    tag_regs1_23 = 54'h0;
  end
  if (reset) begin
    tag_regs1_24 = 54'h0;
  end
  if (reset) begin
    tag_regs1_25 = 54'h0;
  end
  if (reset) begin
    tag_regs1_26 = 54'h0;
  end
  if (reset) begin
    tag_regs1_27 = 54'h0;
  end
  if (reset) begin
    tag_regs1_28 = 54'h0;
  end
  if (reset) begin
    tag_regs1_29 = 54'h0;
  end
  if (reset) begin
    tag_regs1_30 = 54'h0;
  end
  if (reset) begin
    tag_regs1_31 = 54'h0;
  end
  if (reset) begin
    tag_regs1_32 = 54'h0;
  end
  if (reset) begin
    tag_regs1_33 = 54'h0;
  end
  if (reset) begin
    tag_regs1_34 = 54'h0;
  end
  if (reset) begin
    tag_regs1_35 = 54'h0;
  end
  if (reset) begin
    tag_regs1_36 = 54'h0;
  end
  if (reset) begin
    tag_regs1_37 = 54'h0;
  end
  if (reset) begin
    tag_regs1_38 = 54'h0;
  end
  if (reset) begin
    tag_regs1_39 = 54'h0;
  end
  if (reset) begin
    tag_regs1_40 = 54'h0;
  end
  if (reset) begin
    tag_regs1_41 = 54'h0;
  end
  if (reset) begin
    tag_regs1_42 = 54'h0;
  end
  if (reset) begin
    tag_regs1_43 = 54'h0;
  end
  if (reset) begin
    tag_regs1_44 = 54'h0;
  end
  if (reset) begin
    tag_regs1_45 = 54'h0;
  end
  if (reset) begin
    tag_regs1_46 = 54'h0;
  end
  if (reset) begin
    tag_regs1_47 = 54'h0;
  end
  if (reset) begin
    tag_regs1_48 = 54'h0;
  end
  if (reset) begin
    tag_regs1_49 = 54'h0;
  end
  if (reset) begin
    tag_regs1_50 = 54'h0;
  end
  if (reset) begin
    tag_regs1_51 = 54'h0;
  end
  if (reset) begin
    tag_regs1_52 = 54'h0;
  end
  if (reset) begin
    tag_regs1_53 = 54'h0;
  end
  if (reset) begin
    tag_regs1_54 = 54'h0;
  end
  if (reset) begin
    tag_regs1_55 = 54'h0;
  end
  if (reset) begin
    tag_regs1_56 = 54'h0;
  end
  if (reset) begin
    tag_regs1_57 = 54'h0;
  end
  if (reset) begin
    tag_regs1_58 = 54'h0;
  end
  if (reset) begin
    tag_regs1_59 = 54'h0;
  end
  if (reset) begin
    tag_regs1_60 = 54'h0;
  end
  if (reset) begin
    tag_regs1_61 = 54'h0;
  end
  if (reset) begin
    tag_regs1_62 = 54'h0;
  end
  if (reset) begin
    tag_regs1_63 = 54'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module dcache_data(
  input         clock,
  input  [7:0]  io_wen,
  input  [63:0] io_addr,
  input  [63:0] io_wdata,
  output [63:0] io_rdata
);
  wire  dcache_data_ram_0_clock; // @[dcache_data.scala 33:35]
  wire [7:0] dcache_data_ram_0_io_wea; // @[dcache_data.scala 33:35]
  wire [6:0] dcache_data_ram_0_io_addra; // @[dcache_data.scala 33:35]
  wire [63:0] dcache_data_ram_0_io_dina; // @[dcache_data.scala 33:35]
  wire [63:0] dcache_data_ram_0_io_douta; // @[dcache_data.scala 33:35]
  ysyx_sram_with_mask dcache_data_ram_0 ( // @[dcache_data.scala 33:35]
    .clock(dcache_data_ram_0_clock),
    .io_wea(dcache_data_ram_0_io_wea),
    .io_addra(dcache_data_ram_0_io_addra),
    .io_dina(dcache_data_ram_0_io_dina),
    .io_douta(dcache_data_ram_0_io_douta)
  );
  assign io_rdata = dcache_data_ram_0_io_douta; // @[dcache_data.scala 39:16]
  assign dcache_data_ram_0_clock = clock;
  assign dcache_data_ram_0_io_wea = io_wen; // @[dcache_data.scala 35:31]
  assign dcache_data_ram_0_io_addra = io_addr[10:4]; // @[dcache_data.scala 36:42]
  assign dcache_data_ram_0_io_dina = io_wdata; // @[dcache_data.scala 37:31]
endmodule
module data_cache(
  input         clock,
  input         reset,
  output [63:0] io_port_araddr,
  output [3:0]  io_port_arlen,
  output [2:0]  io_port_arsize,
  output [1:0]  io_port_arburst,
  output        io_port_arvalid,
  input         io_port_arready,
  input  [63:0] io_port_rdata,
  input         io_port_rlast,
  input         io_port_rvalid,
  output [63:0] io_port_awaddr,
  output [3:0]  io_port_awlen,
  output [2:0]  io_port_awsize,
  output [1:0]  io_port_awburst,
  output        io_port_awvalid,
  input         io_port_awready,
  output [63:0] io_port_wdata,
  output [7:0]  io_port_wstrb,
  output        io_port_wlast,
  output        io_port_wvalid,
  input         io_port_wready,
  input         io_port_bvalid,
  output        io_stage2_stall,
  output [63:0] io_v_addr_for_tlb,
  input  [63:0] io_p_addr_for_tlb,
  output        io_tlb_req,
  input  [7:0]  io_data_wstrb,
  input         io_sram_req,
  input         io_sram_wr,
  input  [2:0]  io_sram_size,
  input  [63:0] io_sram_addr,
  input  [63:0] io_sram_wdata,
  output [63:0] io_sram_rdata,
  input         io_sram_cache,
  input         io_fence_i_control
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [63:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [63:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [63:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [63:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [63:0] _RAND_406;
  reg [31:0] _RAND_407;
`endif // RANDOMIZE_REG_INIT
  wire  dcache_tag_clock; // @[data_cache.scala 60:30]
  wire  dcache_tag_reset; // @[data_cache.scala 60:30]
  wire  dcache_tag_io_wen; // @[data_cache.scala 60:30]
  wire [53:0] dcache_tag_io_wdata; // @[data_cache.scala 60:30]
  wire [63:0] dcache_tag_io_raddr; // @[data_cache.scala 60:30]
  wire [63:0] dcache_tag_io_waddr; // @[data_cache.scala 60:30]
  wire  dcache_tag_io_hit; // @[data_cache.scala 60:30]
  wire  dcache_tag_io_valid; // @[data_cache.scala 60:30]
  wire [52:0] dcache_tag_io_tag; // @[data_cache.scala 60:30]
  wire  dcache_tag_io_w_valid; // @[data_cache.scala 60:30]
  wire  dcache_tag_1_clock; // @[data_cache.scala 61:30]
  wire  dcache_tag_1_reset; // @[data_cache.scala 61:30]
  wire  dcache_tag_1_io_wen; // @[data_cache.scala 61:30]
  wire [53:0] dcache_tag_1_io_wdata; // @[data_cache.scala 61:30]
  wire [63:0] dcache_tag_1_io_raddr; // @[data_cache.scala 61:30]
  wire [63:0] dcache_tag_1_io_waddr; // @[data_cache.scala 61:30]
  wire  dcache_tag_1_io_hit; // @[data_cache.scala 61:30]
  wire  dcache_tag_1_io_valid; // @[data_cache.scala 61:30]
  wire [52:0] dcache_tag_1_io_tag; // @[data_cache.scala 61:30]
  wire  dcache_tag_1_io_w_valid; // @[data_cache.scala 61:30]
  wire  dcache_data_clock; // @[data_cache.scala 93:62]
  wire [7:0] dcache_data_io_wen; // @[data_cache.scala 93:62]
  wire [63:0] dcache_data_io_addr; // @[data_cache.scala 93:62]
  wire [63:0] dcache_data_io_wdata; // @[data_cache.scala 93:62]
  wire [63:0] dcache_data_io_rdata; // @[data_cache.scala 93:62]
  wire  dcache_data_1_clock; // @[data_cache.scala 93:62]
  wire [7:0] dcache_data_1_io_wen; // @[data_cache.scala 93:62]
  wire [63:0] dcache_data_1_io_addr; // @[data_cache.scala 93:62]
  wire [63:0] dcache_data_1_io_wdata; // @[data_cache.scala 93:62]
  wire [63:0] dcache_data_1_io_rdata; // @[data_cache.scala 93:62]
  wire  dcache_data_2_clock; // @[data_cache.scala 94:62]
  wire [7:0] dcache_data_2_io_wen; // @[data_cache.scala 94:62]
  wire [63:0] dcache_data_2_io_addr; // @[data_cache.scala 94:62]
  wire [63:0] dcache_data_2_io_wdata; // @[data_cache.scala 94:62]
  wire [63:0] dcache_data_2_io_rdata; // @[data_cache.scala 94:62]
  wire  dcache_data_3_clock; // @[data_cache.scala 94:62]
  wire [7:0] dcache_data_3_io_wen; // @[data_cache.scala 94:62]
  wire [63:0] dcache_data_3_io_addr; // @[data_cache.scala 94:62]
  wire [63:0] dcache_data_3_io_wdata; // @[data_cache.scala 94:62]
  wire [63:0] dcache_data_3_io_rdata; // @[data_cache.scala 94:62]
  reg [4:0] work_state; // @[data_cache.scala 53:29]
  reg [2:0] write_counter; // @[data_cache.scala 55:33]
  reg [2:0] read_counter; // @[data_cache.scala 56:32]
  reg [63:0] wait_data; // @[data_cache.scala 57:29]
  reg  lru_0; // @[data_cache.scala 63:22]
  reg  lru_1; // @[data_cache.scala 63:22]
  reg  lru_2; // @[data_cache.scala 63:22]
  reg  lru_3; // @[data_cache.scala 63:22]
  reg  lru_4; // @[data_cache.scala 63:22]
  reg  lru_5; // @[data_cache.scala 63:22]
  reg  lru_6; // @[data_cache.scala 63:22]
  reg  lru_7; // @[data_cache.scala 63:22]
  reg  lru_8; // @[data_cache.scala 63:22]
  reg  lru_9; // @[data_cache.scala 63:22]
  reg  lru_10; // @[data_cache.scala 63:22]
  reg  lru_11; // @[data_cache.scala 63:22]
  reg  lru_12; // @[data_cache.scala 63:22]
  reg  lru_13; // @[data_cache.scala 63:22]
  reg  lru_14; // @[data_cache.scala 63:22]
  reg  lru_15; // @[data_cache.scala 63:22]
  reg  lru_16; // @[data_cache.scala 63:22]
  reg  lru_17; // @[data_cache.scala 63:22]
  reg  lru_18; // @[data_cache.scala 63:22]
  reg  lru_19; // @[data_cache.scala 63:22]
  reg  lru_20; // @[data_cache.scala 63:22]
  reg  lru_21; // @[data_cache.scala 63:22]
  reg  lru_22; // @[data_cache.scala 63:22]
  reg  lru_23; // @[data_cache.scala 63:22]
  reg  lru_24; // @[data_cache.scala 63:22]
  reg  lru_25; // @[data_cache.scala 63:22]
  reg  lru_26; // @[data_cache.scala 63:22]
  reg  lru_27; // @[data_cache.scala 63:22]
  reg  lru_28; // @[data_cache.scala 63:22]
  reg  lru_29; // @[data_cache.scala 63:22]
  reg  lru_30; // @[data_cache.scala 63:22]
  reg  lru_31; // @[data_cache.scala 63:22]
  reg  lru_32; // @[data_cache.scala 63:22]
  reg  lru_33; // @[data_cache.scala 63:22]
  reg  lru_34; // @[data_cache.scala 63:22]
  reg  lru_35; // @[data_cache.scala 63:22]
  reg  lru_36; // @[data_cache.scala 63:22]
  reg  lru_37; // @[data_cache.scala 63:22]
  reg  lru_38; // @[data_cache.scala 63:22]
  reg  lru_39; // @[data_cache.scala 63:22]
  reg  lru_40; // @[data_cache.scala 63:22]
  reg  lru_41; // @[data_cache.scala 63:22]
  reg  lru_42; // @[data_cache.scala 63:22]
  reg  lru_43; // @[data_cache.scala 63:22]
  reg  lru_44; // @[data_cache.scala 63:22]
  reg  lru_45; // @[data_cache.scala 63:22]
  reg  lru_46; // @[data_cache.scala 63:22]
  reg  lru_47; // @[data_cache.scala 63:22]
  reg  lru_48; // @[data_cache.scala 63:22]
  reg  lru_49; // @[data_cache.scala 63:22]
  reg  lru_50; // @[data_cache.scala 63:22]
  reg  lru_51; // @[data_cache.scala 63:22]
  reg  lru_52; // @[data_cache.scala 63:22]
  reg  lru_53; // @[data_cache.scala 63:22]
  reg  lru_54; // @[data_cache.scala 63:22]
  reg  lru_55; // @[data_cache.scala 63:22]
  reg  lru_56; // @[data_cache.scala 63:22]
  reg  lru_57; // @[data_cache.scala 63:22]
  reg  lru_58; // @[data_cache.scala 63:22]
  reg  lru_59; // @[data_cache.scala 63:22]
  reg  lru_60; // @[data_cache.scala 63:22]
  reg  lru_61; // @[data_cache.scala 63:22]
  reg  lru_62; // @[data_cache.scala 63:22]
  reg  lru_63; // @[data_cache.scala 63:22]
  reg  lru_64; // @[data_cache.scala 63:22]
  reg  lru_65; // @[data_cache.scala 63:22]
  reg  lru_66; // @[data_cache.scala 63:22]
  reg  lru_67; // @[data_cache.scala 63:22]
  reg  lru_68; // @[data_cache.scala 63:22]
  reg  lru_69; // @[data_cache.scala 63:22]
  reg  lru_70; // @[data_cache.scala 63:22]
  reg  lru_71; // @[data_cache.scala 63:22]
  reg  lru_72; // @[data_cache.scala 63:22]
  reg  lru_73; // @[data_cache.scala 63:22]
  reg  lru_74; // @[data_cache.scala 63:22]
  reg  lru_75; // @[data_cache.scala 63:22]
  reg  lru_76; // @[data_cache.scala 63:22]
  reg  lru_77; // @[data_cache.scala 63:22]
  reg  lru_78; // @[data_cache.scala 63:22]
  reg  lru_79; // @[data_cache.scala 63:22]
  reg  lru_80; // @[data_cache.scala 63:22]
  reg  lru_81; // @[data_cache.scala 63:22]
  reg  lru_82; // @[data_cache.scala 63:22]
  reg  lru_83; // @[data_cache.scala 63:22]
  reg  lru_84; // @[data_cache.scala 63:22]
  reg  lru_85; // @[data_cache.scala 63:22]
  reg  lru_86; // @[data_cache.scala 63:22]
  reg  lru_87; // @[data_cache.scala 63:22]
  reg  lru_88; // @[data_cache.scala 63:22]
  reg  lru_89; // @[data_cache.scala 63:22]
  reg  lru_90; // @[data_cache.scala 63:22]
  reg  lru_91; // @[data_cache.scala 63:22]
  reg  lru_92; // @[data_cache.scala 63:22]
  reg  lru_93; // @[data_cache.scala 63:22]
  reg  lru_94; // @[data_cache.scala 63:22]
  reg  lru_95; // @[data_cache.scala 63:22]
  reg  lru_96; // @[data_cache.scala 63:22]
  reg  lru_97; // @[data_cache.scala 63:22]
  reg  lru_98; // @[data_cache.scala 63:22]
  reg  lru_99; // @[data_cache.scala 63:22]
  reg  lru_100; // @[data_cache.scala 63:22]
  reg  lru_101; // @[data_cache.scala 63:22]
  reg  lru_102; // @[data_cache.scala 63:22]
  reg  lru_103; // @[data_cache.scala 63:22]
  reg  lru_104; // @[data_cache.scala 63:22]
  reg  lru_105; // @[data_cache.scala 63:22]
  reg  lru_106; // @[data_cache.scala 63:22]
  reg  lru_107; // @[data_cache.scala 63:22]
  reg  lru_108; // @[data_cache.scala 63:22]
  reg  lru_109; // @[data_cache.scala 63:22]
  reg  lru_110; // @[data_cache.scala 63:22]
  reg  lru_111; // @[data_cache.scala 63:22]
  reg  lru_112; // @[data_cache.scala 63:22]
  reg  lru_113; // @[data_cache.scala 63:22]
  reg  lru_114; // @[data_cache.scala 63:22]
  reg  lru_115; // @[data_cache.scala 63:22]
  reg  lru_116; // @[data_cache.scala 63:22]
  reg  lru_117; // @[data_cache.scala 63:22]
  reg  lru_118; // @[data_cache.scala 63:22]
  reg  lru_119; // @[data_cache.scala 63:22]
  reg  lru_120; // @[data_cache.scala 63:22]
  reg  lru_121; // @[data_cache.scala 63:22]
  reg  lru_122; // @[data_cache.scala 63:22]
  reg  lru_123; // @[data_cache.scala 63:22]
  reg  lru_124; // @[data_cache.scala 63:22]
  reg  lru_125; // @[data_cache.scala 63:22]
  reg  lru_126; // @[data_cache.scala 63:22]
  reg  lru_127; // @[data_cache.scala 63:22]
  reg  way0_dirty_0; // @[data_cache.scala 64:29]
  reg  way0_dirty_1; // @[data_cache.scala 64:29]
  reg  way0_dirty_2; // @[data_cache.scala 64:29]
  reg  way0_dirty_3; // @[data_cache.scala 64:29]
  reg  way0_dirty_4; // @[data_cache.scala 64:29]
  reg  way0_dirty_5; // @[data_cache.scala 64:29]
  reg  way0_dirty_6; // @[data_cache.scala 64:29]
  reg  way0_dirty_7; // @[data_cache.scala 64:29]
  reg  way0_dirty_8; // @[data_cache.scala 64:29]
  reg  way0_dirty_9; // @[data_cache.scala 64:29]
  reg  way0_dirty_10; // @[data_cache.scala 64:29]
  reg  way0_dirty_11; // @[data_cache.scala 64:29]
  reg  way0_dirty_12; // @[data_cache.scala 64:29]
  reg  way0_dirty_13; // @[data_cache.scala 64:29]
  reg  way0_dirty_14; // @[data_cache.scala 64:29]
  reg  way0_dirty_15; // @[data_cache.scala 64:29]
  reg  way0_dirty_16; // @[data_cache.scala 64:29]
  reg  way0_dirty_17; // @[data_cache.scala 64:29]
  reg  way0_dirty_18; // @[data_cache.scala 64:29]
  reg  way0_dirty_19; // @[data_cache.scala 64:29]
  reg  way0_dirty_20; // @[data_cache.scala 64:29]
  reg  way0_dirty_21; // @[data_cache.scala 64:29]
  reg  way0_dirty_22; // @[data_cache.scala 64:29]
  reg  way0_dirty_23; // @[data_cache.scala 64:29]
  reg  way0_dirty_24; // @[data_cache.scala 64:29]
  reg  way0_dirty_25; // @[data_cache.scala 64:29]
  reg  way0_dirty_26; // @[data_cache.scala 64:29]
  reg  way0_dirty_27; // @[data_cache.scala 64:29]
  reg  way0_dirty_28; // @[data_cache.scala 64:29]
  reg  way0_dirty_29; // @[data_cache.scala 64:29]
  reg  way0_dirty_30; // @[data_cache.scala 64:29]
  reg  way0_dirty_31; // @[data_cache.scala 64:29]
  reg  way0_dirty_32; // @[data_cache.scala 64:29]
  reg  way0_dirty_33; // @[data_cache.scala 64:29]
  reg  way0_dirty_34; // @[data_cache.scala 64:29]
  reg  way0_dirty_35; // @[data_cache.scala 64:29]
  reg  way0_dirty_36; // @[data_cache.scala 64:29]
  reg  way0_dirty_37; // @[data_cache.scala 64:29]
  reg  way0_dirty_38; // @[data_cache.scala 64:29]
  reg  way0_dirty_39; // @[data_cache.scala 64:29]
  reg  way0_dirty_40; // @[data_cache.scala 64:29]
  reg  way0_dirty_41; // @[data_cache.scala 64:29]
  reg  way0_dirty_42; // @[data_cache.scala 64:29]
  reg  way0_dirty_43; // @[data_cache.scala 64:29]
  reg  way0_dirty_44; // @[data_cache.scala 64:29]
  reg  way0_dirty_45; // @[data_cache.scala 64:29]
  reg  way0_dirty_46; // @[data_cache.scala 64:29]
  reg  way0_dirty_47; // @[data_cache.scala 64:29]
  reg  way0_dirty_48; // @[data_cache.scala 64:29]
  reg  way0_dirty_49; // @[data_cache.scala 64:29]
  reg  way0_dirty_50; // @[data_cache.scala 64:29]
  reg  way0_dirty_51; // @[data_cache.scala 64:29]
  reg  way0_dirty_52; // @[data_cache.scala 64:29]
  reg  way0_dirty_53; // @[data_cache.scala 64:29]
  reg  way0_dirty_54; // @[data_cache.scala 64:29]
  reg  way0_dirty_55; // @[data_cache.scala 64:29]
  reg  way0_dirty_56; // @[data_cache.scala 64:29]
  reg  way0_dirty_57; // @[data_cache.scala 64:29]
  reg  way0_dirty_58; // @[data_cache.scala 64:29]
  reg  way0_dirty_59; // @[data_cache.scala 64:29]
  reg  way0_dirty_60; // @[data_cache.scala 64:29]
  reg  way0_dirty_61; // @[data_cache.scala 64:29]
  reg  way0_dirty_62; // @[data_cache.scala 64:29]
  reg  way0_dirty_63; // @[data_cache.scala 64:29]
  reg  way0_dirty_64; // @[data_cache.scala 64:29]
  reg  way0_dirty_65; // @[data_cache.scala 64:29]
  reg  way0_dirty_66; // @[data_cache.scala 64:29]
  reg  way0_dirty_67; // @[data_cache.scala 64:29]
  reg  way0_dirty_68; // @[data_cache.scala 64:29]
  reg  way0_dirty_69; // @[data_cache.scala 64:29]
  reg  way0_dirty_70; // @[data_cache.scala 64:29]
  reg  way0_dirty_71; // @[data_cache.scala 64:29]
  reg  way0_dirty_72; // @[data_cache.scala 64:29]
  reg  way0_dirty_73; // @[data_cache.scala 64:29]
  reg  way0_dirty_74; // @[data_cache.scala 64:29]
  reg  way0_dirty_75; // @[data_cache.scala 64:29]
  reg  way0_dirty_76; // @[data_cache.scala 64:29]
  reg  way0_dirty_77; // @[data_cache.scala 64:29]
  reg  way0_dirty_78; // @[data_cache.scala 64:29]
  reg  way0_dirty_79; // @[data_cache.scala 64:29]
  reg  way0_dirty_80; // @[data_cache.scala 64:29]
  reg  way0_dirty_81; // @[data_cache.scala 64:29]
  reg  way0_dirty_82; // @[data_cache.scala 64:29]
  reg  way0_dirty_83; // @[data_cache.scala 64:29]
  reg  way0_dirty_84; // @[data_cache.scala 64:29]
  reg  way0_dirty_85; // @[data_cache.scala 64:29]
  reg  way0_dirty_86; // @[data_cache.scala 64:29]
  reg  way0_dirty_87; // @[data_cache.scala 64:29]
  reg  way0_dirty_88; // @[data_cache.scala 64:29]
  reg  way0_dirty_89; // @[data_cache.scala 64:29]
  reg  way0_dirty_90; // @[data_cache.scala 64:29]
  reg  way0_dirty_91; // @[data_cache.scala 64:29]
  reg  way0_dirty_92; // @[data_cache.scala 64:29]
  reg  way0_dirty_93; // @[data_cache.scala 64:29]
  reg  way0_dirty_94; // @[data_cache.scala 64:29]
  reg  way0_dirty_95; // @[data_cache.scala 64:29]
  reg  way0_dirty_96; // @[data_cache.scala 64:29]
  reg  way0_dirty_97; // @[data_cache.scala 64:29]
  reg  way0_dirty_98; // @[data_cache.scala 64:29]
  reg  way0_dirty_99; // @[data_cache.scala 64:29]
  reg  way0_dirty_100; // @[data_cache.scala 64:29]
  reg  way0_dirty_101; // @[data_cache.scala 64:29]
  reg  way0_dirty_102; // @[data_cache.scala 64:29]
  reg  way0_dirty_103; // @[data_cache.scala 64:29]
  reg  way0_dirty_104; // @[data_cache.scala 64:29]
  reg  way0_dirty_105; // @[data_cache.scala 64:29]
  reg  way0_dirty_106; // @[data_cache.scala 64:29]
  reg  way0_dirty_107; // @[data_cache.scala 64:29]
  reg  way0_dirty_108; // @[data_cache.scala 64:29]
  reg  way0_dirty_109; // @[data_cache.scala 64:29]
  reg  way0_dirty_110; // @[data_cache.scala 64:29]
  reg  way0_dirty_111; // @[data_cache.scala 64:29]
  reg  way0_dirty_112; // @[data_cache.scala 64:29]
  reg  way0_dirty_113; // @[data_cache.scala 64:29]
  reg  way0_dirty_114; // @[data_cache.scala 64:29]
  reg  way0_dirty_115; // @[data_cache.scala 64:29]
  reg  way0_dirty_116; // @[data_cache.scala 64:29]
  reg  way0_dirty_117; // @[data_cache.scala 64:29]
  reg  way0_dirty_118; // @[data_cache.scala 64:29]
  reg  way0_dirty_119; // @[data_cache.scala 64:29]
  reg  way0_dirty_120; // @[data_cache.scala 64:29]
  reg  way0_dirty_121; // @[data_cache.scala 64:29]
  reg  way0_dirty_122; // @[data_cache.scala 64:29]
  reg  way0_dirty_123; // @[data_cache.scala 64:29]
  reg  way0_dirty_124; // @[data_cache.scala 64:29]
  reg  way0_dirty_125; // @[data_cache.scala 64:29]
  reg  way0_dirty_126; // @[data_cache.scala 64:29]
  reg  way0_dirty_127; // @[data_cache.scala 64:29]
  reg  way1_dirty_0; // @[data_cache.scala 65:29]
  reg  way1_dirty_1; // @[data_cache.scala 65:29]
  reg  way1_dirty_2; // @[data_cache.scala 65:29]
  reg  way1_dirty_3; // @[data_cache.scala 65:29]
  reg  way1_dirty_4; // @[data_cache.scala 65:29]
  reg  way1_dirty_5; // @[data_cache.scala 65:29]
  reg  way1_dirty_6; // @[data_cache.scala 65:29]
  reg  way1_dirty_7; // @[data_cache.scala 65:29]
  reg  way1_dirty_8; // @[data_cache.scala 65:29]
  reg  way1_dirty_9; // @[data_cache.scala 65:29]
  reg  way1_dirty_10; // @[data_cache.scala 65:29]
  reg  way1_dirty_11; // @[data_cache.scala 65:29]
  reg  way1_dirty_12; // @[data_cache.scala 65:29]
  reg  way1_dirty_13; // @[data_cache.scala 65:29]
  reg  way1_dirty_14; // @[data_cache.scala 65:29]
  reg  way1_dirty_15; // @[data_cache.scala 65:29]
  reg  way1_dirty_16; // @[data_cache.scala 65:29]
  reg  way1_dirty_17; // @[data_cache.scala 65:29]
  reg  way1_dirty_18; // @[data_cache.scala 65:29]
  reg  way1_dirty_19; // @[data_cache.scala 65:29]
  reg  way1_dirty_20; // @[data_cache.scala 65:29]
  reg  way1_dirty_21; // @[data_cache.scala 65:29]
  reg  way1_dirty_22; // @[data_cache.scala 65:29]
  reg  way1_dirty_23; // @[data_cache.scala 65:29]
  reg  way1_dirty_24; // @[data_cache.scala 65:29]
  reg  way1_dirty_25; // @[data_cache.scala 65:29]
  reg  way1_dirty_26; // @[data_cache.scala 65:29]
  reg  way1_dirty_27; // @[data_cache.scala 65:29]
  reg  way1_dirty_28; // @[data_cache.scala 65:29]
  reg  way1_dirty_29; // @[data_cache.scala 65:29]
  reg  way1_dirty_30; // @[data_cache.scala 65:29]
  reg  way1_dirty_31; // @[data_cache.scala 65:29]
  reg  way1_dirty_32; // @[data_cache.scala 65:29]
  reg  way1_dirty_33; // @[data_cache.scala 65:29]
  reg  way1_dirty_34; // @[data_cache.scala 65:29]
  reg  way1_dirty_35; // @[data_cache.scala 65:29]
  reg  way1_dirty_36; // @[data_cache.scala 65:29]
  reg  way1_dirty_37; // @[data_cache.scala 65:29]
  reg  way1_dirty_38; // @[data_cache.scala 65:29]
  reg  way1_dirty_39; // @[data_cache.scala 65:29]
  reg  way1_dirty_40; // @[data_cache.scala 65:29]
  reg  way1_dirty_41; // @[data_cache.scala 65:29]
  reg  way1_dirty_42; // @[data_cache.scala 65:29]
  reg  way1_dirty_43; // @[data_cache.scala 65:29]
  reg  way1_dirty_44; // @[data_cache.scala 65:29]
  reg  way1_dirty_45; // @[data_cache.scala 65:29]
  reg  way1_dirty_46; // @[data_cache.scala 65:29]
  reg  way1_dirty_47; // @[data_cache.scala 65:29]
  reg  way1_dirty_48; // @[data_cache.scala 65:29]
  reg  way1_dirty_49; // @[data_cache.scala 65:29]
  reg  way1_dirty_50; // @[data_cache.scala 65:29]
  reg  way1_dirty_51; // @[data_cache.scala 65:29]
  reg  way1_dirty_52; // @[data_cache.scala 65:29]
  reg  way1_dirty_53; // @[data_cache.scala 65:29]
  reg  way1_dirty_54; // @[data_cache.scala 65:29]
  reg  way1_dirty_55; // @[data_cache.scala 65:29]
  reg  way1_dirty_56; // @[data_cache.scala 65:29]
  reg  way1_dirty_57; // @[data_cache.scala 65:29]
  reg  way1_dirty_58; // @[data_cache.scala 65:29]
  reg  way1_dirty_59; // @[data_cache.scala 65:29]
  reg  way1_dirty_60; // @[data_cache.scala 65:29]
  reg  way1_dirty_61; // @[data_cache.scala 65:29]
  reg  way1_dirty_62; // @[data_cache.scala 65:29]
  reg  way1_dirty_63; // @[data_cache.scala 65:29]
  reg  way1_dirty_64; // @[data_cache.scala 65:29]
  reg  way1_dirty_65; // @[data_cache.scala 65:29]
  reg  way1_dirty_66; // @[data_cache.scala 65:29]
  reg  way1_dirty_67; // @[data_cache.scala 65:29]
  reg  way1_dirty_68; // @[data_cache.scala 65:29]
  reg  way1_dirty_69; // @[data_cache.scala 65:29]
  reg  way1_dirty_70; // @[data_cache.scala 65:29]
  reg  way1_dirty_71; // @[data_cache.scala 65:29]
  reg  way1_dirty_72; // @[data_cache.scala 65:29]
  reg  way1_dirty_73; // @[data_cache.scala 65:29]
  reg  way1_dirty_74; // @[data_cache.scala 65:29]
  reg  way1_dirty_75; // @[data_cache.scala 65:29]
  reg  way1_dirty_76; // @[data_cache.scala 65:29]
  reg  way1_dirty_77; // @[data_cache.scala 65:29]
  reg  way1_dirty_78; // @[data_cache.scala 65:29]
  reg  way1_dirty_79; // @[data_cache.scala 65:29]
  reg  way1_dirty_80; // @[data_cache.scala 65:29]
  reg  way1_dirty_81; // @[data_cache.scala 65:29]
  reg  way1_dirty_82; // @[data_cache.scala 65:29]
  reg  way1_dirty_83; // @[data_cache.scala 65:29]
  reg  way1_dirty_84; // @[data_cache.scala 65:29]
  reg  way1_dirty_85; // @[data_cache.scala 65:29]
  reg  way1_dirty_86; // @[data_cache.scala 65:29]
  reg  way1_dirty_87; // @[data_cache.scala 65:29]
  reg  way1_dirty_88; // @[data_cache.scala 65:29]
  reg  way1_dirty_89; // @[data_cache.scala 65:29]
  reg  way1_dirty_90; // @[data_cache.scala 65:29]
  reg  way1_dirty_91; // @[data_cache.scala 65:29]
  reg  way1_dirty_92; // @[data_cache.scala 65:29]
  reg  way1_dirty_93; // @[data_cache.scala 65:29]
  reg  way1_dirty_94; // @[data_cache.scala 65:29]
  reg  way1_dirty_95; // @[data_cache.scala 65:29]
  reg  way1_dirty_96; // @[data_cache.scala 65:29]
  reg  way1_dirty_97; // @[data_cache.scala 65:29]
  reg  way1_dirty_98; // @[data_cache.scala 65:29]
  reg  way1_dirty_99; // @[data_cache.scala 65:29]
  reg  way1_dirty_100; // @[data_cache.scala 65:29]
  reg  way1_dirty_101; // @[data_cache.scala 65:29]
  reg  way1_dirty_102; // @[data_cache.scala 65:29]
  reg  way1_dirty_103; // @[data_cache.scala 65:29]
  reg  way1_dirty_104; // @[data_cache.scala 65:29]
  reg  way1_dirty_105; // @[data_cache.scala 65:29]
  reg  way1_dirty_106; // @[data_cache.scala 65:29]
  reg  way1_dirty_107; // @[data_cache.scala 65:29]
  reg  way1_dirty_108; // @[data_cache.scala 65:29]
  reg  way1_dirty_109; // @[data_cache.scala 65:29]
  reg  way1_dirty_110; // @[data_cache.scala 65:29]
  reg  way1_dirty_111; // @[data_cache.scala 65:29]
  reg  way1_dirty_112; // @[data_cache.scala 65:29]
  reg  way1_dirty_113; // @[data_cache.scala 65:29]
  reg  way1_dirty_114; // @[data_cache.scala 65:29]
  reg  way1_dirty_115; // @[data_cache.scala 65:29]
  reg  way1_dirty_116; // @[data_cache.scala 65:29]
  reg  way1_dirty_117; // @[data_cache.scala 65:29]
  reg  way1_dirty_118; // @[data_cache.scala 65:29]
  reg  way1_dirty_119; // @[data_cache.scala 65:29]
  reg  way1_dirty_120; // @[data_cache.scala 65:29]
  reg  way1_dirty_121; // @[data_cache.scala 65:29]
  reg  way1_dirty_122; // @[data_cache.scala 65:29]
  reg  way1_dirty_123; // @[data_cache.scala 65:29]
  reg  way1_dirty_124; // @[data_cache.scala 65:29]
  reg  way1_dirty_125; // @[data_cache.scala 65:29]
  reg  way1_dirty_126; // @[data_cache.scala 65:29]
  reg  way1_dirty_127; // @[data_cache.scala 65:29]
  reg [63:0] stage1_addr_line_mapping; // @[data_cache.scala 69:39]
  reg  stage1_sram_cache_reg; // @[data_cache.scala 70:40]
  reg [63:0] stage1_sram_wdata_reg; // @[data_cache.scala 71:40]
  reg [1:0] stage1_sram_size_reg; // @[data_cache.scala 72:39]
  reg  stage1_sram_wr_reg; // @[data_cache.scala 73:37]
  reg  stage1_sram_req_reg; // @[data_cache.scala 74:38]
  reg  stage1_sram_hit0_reg; // @[data_cache.scala 76:40]
  reg  stage1_sram_hit1_reg; // @[data_cache.scala 77:40]
  reg  stage1_sram_valid0_reg; // @[data_cache.scala 78:42]
  reg  stage1_sram_valid1_reg; // @[data_cache.scala 79:42]
  reg [7:0] stage1_wstrb_reg; // @[data_cache.scala 80:35]
  reg [63:0] stage1_sram_phy_addr_reg; // @[data_cache.scala 82:43]
  reg [7:0] data_write_back_counter; // @[data_cache.scala 141:42]
  wire  _data_cache_under_write_back_T = work_state == 5'h11; // @[data_cache.scala 143:51]
  wire  _data_cache_under_write_back_T_1 = work_state == 5'h15; // @[data_cache.scala 143:93]
  wire  _data_cache_under_write_back_T_3 = work_state == 5'h12; // @[data_cache.scala 143:135]
  wire  _data_cache_under_write_back_T_4 = work_state == 5'h11 | work_state == 5'h15 | work_state == 5'h12; // @[data_cache.scala 143:121]
  wire  _data_cache_under_write_back_T_5 = work_state == 5'h13; // @[data_cache.scala 144:23]
  wire  data_cache_under_write_back = _data_cache_under_write_back_T_4 | work_state == 5'h13 | work_state == 5'h14; // @[data_cache.scala 144:53]
  wire  _GEN_1 = 7'h1 == data_write_back_counter[6:0] ? way1_dirty_1 : way1_dirty_0; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_2 = 7'h2 == data_write_back_counter[6:0] ? way1_dirty_2 : _GEN_1; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_3 = 7'h3 == data_write_back_counter[6:0] ? way1_dirty_3 : _GEN_2; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_4 = 7'h4 == data_write_back_counter[6:0] ? way1_dirty_4 : _GEN_3; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_5 = 7'h5 == data_write_back_counter[6:0] ? way1_dirty_5 : _GEN_4; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_6 = 7'h6 == data_write_back_counter[6:0] ? way1_dirty_6 : _GEN_5; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_7 = 7'h7 == data_write_back_counter[6:0] ? way1_dirty_7 : _GEN_6; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_8 = 7'h8 == data_write_back_counter[6:0] ? way1_dirty_8 : _GEN_7; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_9 = 7'h9 == data_write_back_counter[6:0] ? way1_dirty_9 : _GEN_8; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_10 = 7'ha == data_write_back_counter[6:0] ? way1_dirty_10 : _GEN_9; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_11 = 7'hb == data_write_back_counter[6:0] ? way1_dirty_11 : _GEN_10; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_12 = 7'hc == data_write_back_counter[6:0] ? way1_dirty_12 : _GEN_11; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_13 = 7'hd == data_write_back_counter[6:0] ? way1_dirty_13 : _GEN_12; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_14 = 7'he == data_write_back_counter[6:0] ? way1_dirty_14 : _GEN_13; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_15 = 7'hf == data_write_back_counter[6:0] ? way1_dirty_15 : _GEN_14; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_16 = 7'h10 == data_write_back_counter[6:0] ? way1_dirty_16 : _GEN_15; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_17 = 7'h11 == data_write_back_counter[6:0] ? way1_dirty_17 : _GEN_16; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_18 = 7'h12 == data_write_back_counter[6:0] ? way1_dirty_18 : _GEN_17; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_19 = 7'h13 == data_write_back_counter[6:0] ? way1_dirty_19 : _GEN_18; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_20 = 7'h14 == data_write_back_counter[6:0] ? way1_dirty_20 : _GEN_19; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_21 = 7'h15 == data_write_back_counter[6:0] ? way1_dirty_21 : _GEN_20; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_22 = 7'h16 == data_write_back_counter[6:0] ? way1_dirty_22 : _GEN_21; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_23 = 7'h17 == data_write_back_counter[6:0] ? way1_dirty_23 : _GEN_22; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_24 = 7'h18 == data_write_back_counter[6:0] ? way1_dirty_24 : _GEN_23; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_25 = 7'h19 == data_write_back_counter[6:0] ? way1_dirty_25 : _GEN_24; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_26 = 7'h1a == data_write_back_counter[6:0] ? way1_dirty_26 : _GEN_25; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_27 = 7'h1b == data_write_back_counter[6:0] ? way1_dirty_27 : _GEN_26; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_28 = 7'h1c == data_write_back_counter[6:0] ? way1_dirty_28 : _GEN_27; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_29 = 7'h1d == data_write_back_counter[6:0] ? way1_dirty_29 : _GEN_28; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_30 = 7'h1e == data_write_back_counter[6:0] ? way1_dirty_30 : _GEN_29; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_31 = 7'h1f == data_write_back_counter[6:0] ? way1_dirty_31 : _GEN_30; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_32 = 7'h20 == data_write_back_counter[6:0] ? way1_dirty_32 : _GEN_31; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_33 = 7'h21 == data_write_back_counter[6:0] ? way1_dirty_33 : _GEN_32; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_34 = 7'h22 == data_write_back_counter[6:0] ? way1_dirty_34 : _GEN_33; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_35 = 7'h23 == data_write_back_counter[6:0] ? way1_dirty_35 : _GEN_34; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_36 = 7'h24 == data_write_back_counter[6:0] ? way1_dirty_36 : _GEN_35; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_37 = 7'h25 == data_write_back_counter[6:0] ? way1_dirty_37 : _GEN_36; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_38 = 7'h26 == data_write_back_counter[6:0] ? way1_dirty_38 : _GEN_37; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_39 = 7'h27 == data_write_back_counter[6:0] ? way1_dirty_39 : _GEN_38; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_40 = 7'h28 == data_write_back_counter[6:0] ? way1_dirty_40 : _GEN_39; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_41 = 7'h29 == data_write_back_counter[6:0] ? way1_dirty_41 : _GEN_40; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_42 = 7'h2a == data_write_back_counter[6:0] ? way1_dirty_42 : _GEN_41; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_43 = 7'h2b == data_write_back_counter[6:0] ? way1_dirty_43 : _GEN_42; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_44 = 7'h2c == data_write_back_counter[6:0] ? way1_dirty_44 : _GEN_43; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_45 = 7'h2d == data_write_back_counter[6:0] ? way1_dirty_45 : _GEN_44; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_46 = 7'h2e == data_write_back_counter[6:0] ? way1_dirty_46 : _GEN_45; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_47 = 7'h2f == data_write_back_counter[6:0] ? way1_dirty_47 : _GEN_46; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_48 = 7'h30 == data_write_back_counter[6:0] ? way1_dirty_48 : _GEN_47; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_49 = 7'h31 == data_write_back_counter[6:0] ? way1_dirty_49 : _GEN_48; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_50 = 7'h32 == data_write_back_counter[6:0] ? way1_dirty_50 : _GEN_49; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_51 = 7'h33 == data_write_back_counter[6:0] ? way1_dirty_51 : _GEN_50; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_52 = 7'h34 == data_write_back_counter[6:0] ? way1_dirty_52 : _GEN_51; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_53 = 7'h35 == data_write_back_counter[6:0] ? way1_dirty_53 : _GEN_52; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_54 = 7'h36 == data_write_back_counter[6:0] ? way1_dirty_54 : _GEN_53; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_55 = 7'h37 == data_write_back_counter[6:0] ? way1_dirty_55 : _GEN_54; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_56 = 7'h38 == data_write_back_counter[6:0] ? way1_dirty_56 : _GEN_55; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_57 = 7'h39 == data_write_back_counter[6:0] ? way1_dirty_57 : _GEN_56; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_58 = 7'h3a == data_write_back_counter[6:0] ? way1_dirty_58 : _GEN_57; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_59 = 7'h3b == data_write_back_counter[6:0] ? way1_dirty_59 : _GEN_58; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_60 = 7'h3c == data_write_back_counter[6:0] ? way1_dirty_60 : _GEN_59; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_61 = 7'h3d == data_write_back_counter[6:0] ? way1_dirty_61 : _GEN_60; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_62 = 7'h3e == data_write_back_counter[6:0] ? way1_dirty_62 : _GEN_61; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_63 = 7'h3f == data_write_back_counter[6:0] ? way1_dirty_63 : _GEN_62; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_64 = 7'h40 == data_write_back_counter[6:0] ? way1_dirty_64 : _GEN_63; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_65 = 7'h41 == data_write_back_counter[6:0] ? way1_dirty_65 : _GEN_64; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_66 = 7'h42 == data_write_back_counter[6:0] ? way1_dirty_66 : _GEN_65; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_67 = 7'h43 == data_write_back_counter[6:0] ? way1_dirty_67 : _GEN_66; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_68 = 7'h44 == data_write_back_counter[6:0] ? way1_dirty_68 : _GEN_67; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_69 = 7'h45 == data_write_back_counter[6:0] ? way1_dirty_69 : _GEN_68; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_70 = 7'h46 == data_write_back_counter[6:0] ? way1_dirty_70 : _GEN_69; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_71 = 7'h47 == data_write_back_counter[6:0] ? way1_dirty_71 : _GEN_70; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_72 = 7'h48 == data_write_back_counter[6:0] ? way1_dirty_72 : _GEN_71; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_73 = 7'h49 == data_write_back_counter[6:0] ? way1_dirty_73 : _GEN_72; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_74 = 7'h4a == data_write_back_counter[6:0] ? way1_dirty_74 : _GEN_73; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_75 = 7'h4b == data_write_back_counter[6:0] ? way1_dirty_75 : _GEN_74; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_76 = 7'h4c == data_write_back_counter[6:0] ? way1_dirty_76 : _GEN_75; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_77 = 7'h4d == data_write_back_counter[6:0] ? way1_dirty_77 : _GEN_76; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_78 = 7'h4e == data_write_back_counter[6:0] ? way1_dirty_78 : _GEN_77; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_79 = 7'h4f == data_write_back_counter[6:0] ? way1_dirty_79 : _GEN_78; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_80 = 7'h50 == data_write_back_counter[6:0] ? way1_dirty_80 : _GEN_79; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_81 = 7'h51 == data_write_back_counter[6:0] ? way1_dirty_81 : _GEN_80; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_82 = 7'h52 == data_write_back_counter[6:0] ? way1_dirty_82 : _GEN_81; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_83 = 7'h53 == data_write_back_counter[6:0] ? way1_dirty_83 : _GEN_82; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_84 = 7'h54 == data_write_back_counter[6:0] ? way1_dirty_84 : _GEN_83; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_85 = 7'h55 == data_write_back_counter[6:0] ? way1_dirty_85 : _GEN_84; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_86 = 7'h56 == data_write_back_counter[6:0] ? way1_dirty_86 : _GEN_85; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_87 = 7'h57 == data_write_back_counter[6:0] ? way1_dirty_87 : _GEN_86; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_88 = 7'h58 == data_write_back_counter[6:0] ? way1_dirty_88 : _GEN_87; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_89 = 7'h59 == data_write_back_counter[6:0] ? way1_dirty_89 : _GEN_88; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_90 = 7'h5a == data_write_back_counter[6:0] ? way1_dirty_90 : _GEN_89; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_91 = 7'h5b == data_write_back_counter[6:0] ? way1_dirty_91 : _GEN_90; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_92 = 7'h5c == data_write_back_counter[6:0] ? way1_dirty_92 : _GEN_91; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_93 = 7'h5d == data_write_back_counter[6:0] ? way1_dirty_93 : _GEN_92; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_94 = 7'h5e == data_write_back_counter[6:0] ? way1_dirty_94 : _GEN_93; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_95 = 7'h5f == data_write_back_counter[6:0] ? way1_dirty_95 : _GEN_94; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_96 = 7'h60 == data_write_back_counter[6:0] ? way1_dirty_96 : _GEN_95; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_97 = 7'h61 == data_write_back_counter[6:0] ? way1_dirty_97 : _GEN_96; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_98 = 7'h62 == data_write_back_counter[6:0] ? way1_dirty_98 : _GEN_97; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_99 = 7'h63 == data_write_back_counter[6:0] ? way1_dirty_99 : _GEN_98; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_100 = 7'h64 == data_write_back_counter[6:0] ? way1_dirty_100 : _GEN_99; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_101 = 7'h65 == data_write_back_counter[6:0] ? way1_dirty_101 : _GEN_100; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_102 = 7'h66 == data_write_back_counter[6:0] ? way1_dirty_102 : _GEN_101; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_103 = 7'h67 == data_write_back_counter[6:0] ? way1_dirty_103 : _GEN_102; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_104 = 7'h68 == data_write_back_counter[6:0] ? way1_dirty_104 : _GEN_103; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_105 = 7'h69 == data_write_back_counter[6:0] ? way1_dirty_105 : _GEN_104; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_106 = 7'h6a == data_write_back_counter[6:0] ? way1_dirty_106 : _GEN_105; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_107 = 7'h6b == data_write_back_counter[6:0] ? way1_dirty_107 : _GEN_106; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_108 = 7'h6c == data_write_back_counter[6:0] ? way1_dirty_108 : _GEN_107; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_109 = 7'h6d == data_write_back_counter[6:0] ? way1_dirty_109 : _GEN_108; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_110 = 7'h6e == data_write_back_counter[6:0] ? way1_dirty_110 : _GEN_109; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_111 = 7'h6f == data_write_back_counter[6:0] ? way1_dirty_111 : _GEN_110; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_112 = 7'h70 == data_write_back_counter[6:0] ? way1_dirty_112 : _GEN_111; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_113 = 7'h71 == data_write_back_counter[6:0] ? way1_dirty_113 : _GEN_112; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_114 = 7'h72 == data_write_back_counter[6:0] ? way1_dirty_114 : _GEN_113; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_115 = 7'h73 == data_write_back_counter[6:0] ? way1_dirty_115 : _GEN_114; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_116 = 7'h74 == data_write_back_counter[6:0] ? way1_dirty_116 : _GEN_115; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_117 = 7'h75 == data_write_back_counter[6:0] ? way1_dirty_117 : _GEN_116; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_118 = 7'h76 == data_write_back_counter[6:0] ? way1_dirty_118 : _GEN_117; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_119 = 7'h77 == data_write_back_counter[6:0] ? way1_dirty_119 : _GEN_118; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_120 = 7'h78 == data_write_back_counter[6:0] ? way1_dirty_120 : _GEN_119; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_121 = 7'h79 == data_write_back_counter[6:0] ? way1_dirty_121 : _GEN_120; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_122 = 7'h7a == data_write_back_counter[6:0] ? way1_dirty_122 : _GEN_121; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_123 = 7'h7b == data_write_back_counter[6:0] ? way1_dirty_123 : _GEN_122; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_124 = 7'h7c == data_write_back_counter[6:0] ? way1_dirty_124 : _GEN_123; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_125 = 7'h7d == data_write_back_counter[6:0] ? way1_dirty_125 : _GEN_124; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_126 = 7'h7e == data_write_back_counter[6:0] ? way1_dirty_126 : _GEN_125; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_127 = 7'h7f == data_write_back_counter[6:0] ? way1_dirty_127 : _GEN_126; // @[data_cache.scala 154:{149,149}]
  wire  _GEN_129 = 7'h1 == data_write_back_counter[6:0] ? way0_dirty_1 : way0_dirty_0; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_130 = 7'h2 == data_write_back_counter[6:0] ? way0_dirty_2 : _GEN_129; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_131 = 7'h3 == data_write_back_counter[6:0] ? way0_dirty_3 : _GEN_130; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_132 = 7'h4 == data_write_back_counter[6:0] ? way0_dirty_4 : _GEN_131; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_133 = 7'h5 == data_write_back_counter[6:0] ? way0_dirty_5 : _GEN_132; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_134 = 7'h6 == data_write_back_counter[6:0] ? way0_dirty_6 : _GEN_133; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_135 = 7'h7 == data_write_back_counter[6:0] ? way0_dirty_7 : _GEN_134; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_136 = 7'h8 == data_write_back_counter[6:0] ? way0_dirty_8 : _GEN_135; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_137 = 7'h9 == data_write_back_counter[6:0] ? way0_dirty_9 : _GEN_136; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_138 = 7'ha == data_write_back_counter[6:0] ? way0_dirty_10 : _GEN_137; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_139 = 7'hb == data_write_back_counter[6:0] ? way0_dirty_11 : _GEN_138; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_140 = 7'hc == data_write_back_counter[6:0] ? way0_dirty_12 : _GEN_139; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_141 = 7'hd == data_write_back_counter[6:0] ? way0_dirty_13 : _GEN_140; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_142 = 7'he == data_write_back_counter[6:0] ? way0_dirty_14 : _GEN_141; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_143 = 7'hf == data_write_back_counter[6:0] ? way0_dirty_15 : _GEN_142; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_144 = 7'h10 == data_write_back_counter[6:0] ? way0_dirty_16 : _GEN_143; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_145 = 7'h11 == data_write_back_counter[6:0] ? way0_dirty_17 : _GEN_144; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_146 = 7'h12 == data_write_back_counter[6:0] ? way0_dirty_18 : _GEN_145; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_147 = 7'h13 == data_write_back_counter[6:0] ? way0_dirty_19 : _GEN_146; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_148 = 7'h14 == data_write_back_counter[6:0] ? way0_dirty_20 : _GEN_147; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_149 = 7'h15 == data_write_back_counter[6:0] ? way0_dirty_21 : _GEN_148; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_150 = 7'h16 == data_write_back_counter[6:0] ? way0_dirty_22 : _GEN_149; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_151 = 7'h17 == data_write_back_counter[6:0] ? way0_dirty_23 : _GEN_150; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_152 = 7'h18 == data_write_back_counter[6:0] ? way0_dirty_24 : _GEN_151; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_153 = 7'h19 == data_write_back_counter[6:0] ? way0_dirty_25 : _GEN_152; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_154 = 7'h1a == data_write_back_counter[6:0] ? way0_dirty_26 : _GEN_153; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_155 = 7'h1b == data_write_back_counter[6:0] ? way0_dirty_27 : _GEN_154; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_156 = 7'h1c == data_write_back_counter[6:0] ? way0_dirty_28 : _GEN_155; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_157 = 7'h1d == data_write_back_counter[6:0] ? way0_dirty_29 : _GEN_156; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_158 = 7'h1e == data_write_back_counter[6:0] ? way0_dirty_30 : _GEN_157; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_159 = 7'h1f == data_write_back_counter[6:0] ? way0_dirty_31 : _GEN_158; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_160 = 7'h20 == data_write_back_counter[6:0] ? way0_dirty_32 : _GEN_159; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_161 = 7'h21 == data_write_back_counter[6:0] ? way0_dirty_33 : _GEN_160; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_162 = 7'h22 == data_write_back_counter[6:0] ? way0_dirty_34 : _GEN_161; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_163 = 7'h23 == data_write_back_counter[6:0] ? way0_dirty_35 : _GEN_162; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_164 = 7'h24 == data_write_back_counter[6:0] ? way0_dirty_36 : _GEN_163; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_165 = 7'h25 == data_write_back_counter[6:0] ? way0_dirty_37 : _GEN_164; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_166 = 7'h26 == data_write_back_counter[6:0] ? way0_dirty_38 : _GEN_165; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_167 = 7'h27 == data_write_back_counter[6:0] ? way0_dirty_39 : _GEN_166; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_168 = 7'h28 == data_write_back_counter[6:0] ? way0_dirty_40 : _GEN_167; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_169 = 7'h29 == data_write_back_counter[6:0] ? way0_dirty_41 : _GEN_168; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_170 = 7'h2a == data_write_back_counter[6:0] ? way0_dirty_42 : _GEN_169; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_171 = 7'h2b == data_write_back_counter[6:0] ? way0_dirty_43 : _GEN_170; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_172 = 7'h2c == data_write_back_counter[6:0] ? way0_dirty_44 : _GEN_171; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_173 = 7'h2d == data_write_back_counter[6:0] ? way0_dirty_45 : _GEN_172; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_174 = 7'h2e == data_write_back_counter[6:0] ? way0_dirty_46 : _GEN_173; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_175 = 7'h2f == data_write_back_counter[6:0] ? way0_dirty_47 : _GEN_174; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_176 = 7'h30 == data_write_back_counter[6:0] ? way0_dirty_48 : _GEN_175; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_177 = 7'h31 == data_write_back_counter[6:0] ? way0_dirty_49 : _GEN_176; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_178 = 7'h32 == data_write_back_counter[6:0] ? way0_dirty_50 : _GEN_177; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_179 = 7'h33 == data_write_back_counter[6:0] ? way0_dirty_51 : _GEN_178; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_180 = 7'h34 == data_write_back_counter[6:0] ? way0_dirty_52 : _GEN_179; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_181 = 7'h35 == data_write_back_counter[6:0] ? way0_dirty_53 : _GEN_180; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_182 = 7'h36 == data_write_back_counter[6:0] ? way0_dirty_54 : _GEN_181; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_183 = 7'h37 == data_write_back_counter[6:0] ? way0_dirty_55 : _GEN_182; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_184 = 7'h38 == data_write_back_counter[6:0] ? way0_dirty_56 : _GEN_183; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_185 = 7'h39 == data_write_back_counter[6:0] ? way0_dirty_57 : _GEN_184; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_186 = 7'h3a == data_write_back_counter[6:0] ? way0_dirty_58 : _GEN_185; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_187 = 7'h3b == data_write_back_counter[6:0] ? way0_dirty_59 : _GEN_186; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_188 = 7'h3c == data_write_back_counter[6:0] ? way0_dirty_60 : _GEN_187; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_189 = 7'h3d == data_write_back_counter[6:0] ? way0_dirty_61 : _GEN_188; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_190 = 7'h3e == data_write_back_counter[6:0] ? way0_dirty_62 : _GEN_189; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_191 = 7'h3f == data_write_back_counter[6:0] ? way0_dirty_63 : _GEN_190; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_192 = 7'h40 == data_write_back_counter[6:0] ? way0_dirty_64 : _GEN_191; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_193 = 7'h41 == data_write_back_counter[6:0] ? way0_dirty_65 : _GEN_192; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_194 = 7'h42 == data_write_back_counter[6:0] ? way0_dirty_66 : _GEN_193; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_195 = 7'h43 == data_write_back_counter[6:0] ? way0_dirty_67 : _GEN_194; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_196 = 7'h44 == data_write_back_counter[6:0] ? way0_dirty_68 : _GEN_195; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_197 = 7'h45 == data_write_back_counter[6:0] ? way0_dirty_69 : _GEN_196; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_198 = 7'h46 == data_write_back_counter[6:0] ? way0_dirty_70 : _GEN_197; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_199 = 7'h47 == data_write_back_counter[6:0] ? way0_dirty_71 : _GEN_198; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_200 = 7'h48 == data_write_back_counter[6:0] ? way0_dirty_72 : _GEN_199; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_201 = 7'h49 == data_write_back_counter[6:0] ? way0_dirty_73 : _GEN_200; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_202 = 7'h4a == data_write_back_counter[6:0] ? way0_dirty_74 : _GEN_201; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_203 = 7'h4b == data_write_back_counter[6:0] ? way0_dirty_75 : _GEN_202; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_204 = 7'h4c == data_write_back_counter[6:0] ? way0_dirty_76 : _GEN_203; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_205 = 7'h4d == data_write_back_counter[6:0] ? way0_dirty_77 : _GEN_204; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_206 = 7'h4e == data_write_back_counter[6:0] ? way0_dirty_78 : _GEN_205; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_207 = 7'h4f == data_write_back_counter[6:0] ? way0_dirty_79 : _GEN_206; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_208 = 7'h50 == data_write_back_counter[6:0] ? way0_dirty_80 : _GEN_207; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_209 = 7'h51 == data_write_back_counter[6:0] ? way0_dirty_81 : _GEN_208; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_210 = 7'h52 == data_write_back_counter[6:0] ? way0_dirty_82 : _GEN_209; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_211 = 7'h53 == data_write_back_counter[6:0] ? way0_dirty_83 : _GEN_210; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_212 = 7'h54 == data_write_back_counter[6:0] ? way0_dirty_84 : _GEN_211; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_213 = 7'h55 == data_write_back_counter[6:0] ? way0_dirty_85 : _GEN_212; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_214 = 7'h56 == data_write_back_counter[6:0] ? way0_dirty_86 : _GEN_213; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_215 = 7'h57 == data_write_back_counter[6:0] ? way0_dirty_87 : _GEN_214; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_216 = 7'h58 == data_write_back_counter[6:0] ? way0_dirty_88 : _GEN_215; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_217 = 7'h59 == data_write_back_counter[6:0] ? way0_dirty_89 : _GEN_216; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_218 = 7'h5a == data_write_back_counter[6:0] ? way0_dirty_90 : _GEN_217; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_219 = 7'h5b == data_write_back_counter[6:0] ? way0_dirty_91 : _GEN_218; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_220 = 7'h5c == data_write_back_counter[6:0] ? way0_dirty_92 : _GEN_219; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_221 = 7'h5d == data_write_back_counter[6:0] ? way0_dirty_93 : _GEN_220; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_222 = 7'h5e == data_write_back_counter[6:0] ? way0_dirty_94 : _GEN_221; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_223 = 7'h5f == data_write_back_counter[6:0] ? way0_dirty_95 : _GEN_222; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_224 = 7'h60 == data_write_back_counter[6:0] ? way0_dirty_96 : _GEN_223; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_225 = 7'h61 == data_write_back_counter[6:0] ? way0_dirty_97 : _GEN_224; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_226 = 7'h62 == data_write_back_counter[6:0] ? way0_dirty_98 : _GEN_225; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_227 = 7'h63 == data_write_back_counter[6:0] ? way0_dirty_99 : _GEN_226; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_228 = 7'h64 == data_write_back_counter[6:0] ? way0_dirty_100 : _GEN_227; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_229 = 7'h65 == data_write_back_counter[6:0] ? way0_dirty_101 : _GEN_228; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_230 = 7'h66 == data_write_back_counter[6:0] ? way0_dirty_102 : _GEN_229; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_231 = 7'h67 == data_write_back_counter[6:0] ? way0_dirty_103 : _GEN_230; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_232 = 7'h68 == data_write_back_counter[6:0] ? way0_dirty_104 : _GEN_231; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_233 = 7'h69 == data_write_back_counter[6:0] ? way0_dirty_105 : _GEN_232; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_234 = 7'h6a == data_write_back_counter[6:0] ? way0_dirty_106 : _GEN_233; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_235 = 7'h6b == data_write_back_counter[6:0] ? way0_dirty_107 : _GEN_234; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_236 = 7'h6c == data_write_back_counter[6:0] ? way0_dirty_108 : _GEN_235; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_237 = 7'h6d == data_write_back_counter[6:0] ? way0_dirty_109 : _GEN_236; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_238 = 7'h6e == data_write_back_counter[6:0] ? way0_dirty_110 : _GEN_237; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_239 = 7'h6f == data_write_back_counter[6:0] ? way0_dirty_111 : _GEN_238; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_240 = 7'h70 == data_write_back_counter[6:0] ? way0_dirty_112 : _GEN_239; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_241 = 7'h71 == data_write_back_counter[6:0] ? way0_dirty_113 : _GEN_240; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_242 = 7'h72 == data_write_back_counter[6:0] ? way0_dirty_114 : _GEN_241; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_243 = 7'h73 == data_write_back_counter[6:0] ? way0_dirty_115 : _GEN_242; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_244 = 7'h74 == data_write_back_counter[6:0] ? way0_dirty_116 : _GEN_243; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_245 = 7'h75 == data_write_back_counter[6:0] ? way0_dirty_117 : _GEN_244; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_246 = 7'h76 == data_write_back_counter[6:0] ? way0_dirty_118 : _GEN_245; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_247 = 7'h77 == data_write_back_counter[6:0] ? way0_dirty_119 : _GEN_246; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_248 = 7'h78 == data_write_back_counter[6:0] ? way0_dirty_120 : _GEN_247; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_249 = 7'h79 == data_write_back_counter[6:0] ? way0_dirty_121 : _GEN_248; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_250 = 7'h7a == data_write_back_counter[6:0] ? way0_dirty_122 : _GEN_249; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_251 = 7'h7b == data_write_back_counter[6:0] ? way0_dirty_123 : _GEN_250; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_252 = 7'h7c == data_write_back_counter[6:0] ? way0_dirty_124 : _GEN_251; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_253 = 7'h7d == data_write_back_counter[6:0] ? way0_dirty_125 : _GEN_252; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_254 = 7'h7e == data_write_back_counter[6:0] ? way0_dirty_126 : _GEN_253; // @[data_cache.scala 155:{87,87}]
  wire  _GEN_255 = 7'h7f == data_write_back_counter[6:0] ? way0_dirty_127 : _GEN_254; // @[data_cache.scala 155:{87,87}]
  wire  _data_should_write_back_T_6 = dcache_tag_io_w_valid & _GEN_255; // @[data_cache.scala 155:30]
  wire  data_should_write_back = data_write_back_counter[7] ? dcache_tag_1_io_w_valid & _GEN_127 :
    _data_should_write_back_T_6; // @[data_cache.scala 154:34]
  wire  _data_write_back_counter_T_2 = _data_cache_under_write_back_T & ~data_should_write_back; // @[data_cache.scala 148:49]
  wire [7:0] _data_write_back_counter_T_4 = data_write_back_counter + 8'h1; // @[data_cache.scala 148:106]
  wire  data_all_write_back = data_write_back_counter == 8'hff; // @[data_cache.scala 153:55]
  wire  _hit_T = stage1_sram_hit0_reg & stage1_sram_valid0_reg; // @[data_cache.scala 233:37]
  wire  _hit_T_1 = stage1_sram_hit1_reg & stage1_sram_valid1_reg; // @[data_cache.scala 234:31]
  wire  hit = stage1_sram_hit0_reg & stage1_sram_valid0_reg | _hit_T_1; // @[data_cache.scala 233:64]
  wire [4:0] _state_ready_lookup_should_be_T_2 = stage1_sram_cache_reg ? 5'h19 : 5'h0; // @[data_cache.scala 244:82]
  wire [4:0] _state_ready_lookup_should_be_T_3 = stage1_sram_req_reg ? _state_ready_lookup_should_be_T_2 : 5'h19; // @[data_cache.scala 244:51]
  wire [4:0] _state_ready_lookup_should_be_T_5 = stage1_sram_req_reg ? 5'h0 : 5'h19; // @[data_cache.scala 245:16]
  wire [4:0] state_ready_lookup_should_be = hit ? _state_ready_lookup_should_be_T_3 : _state_ready_lookup_should_be_T_5; // @[data_cache.scala 244:43]
  wire [4:0] _access_work_state_for_stall_T_3 = io_port_bvalid ? 5'h18 : 5'h5; // @[data_cache.scala 279:40]
  wire [4:0] _access_work_state_for_stall_T_1 = io_port_rvalid ? 5'h18 : work_state; // @[data_cache.scala 277:39]
  wire [4:0] _access_work_state_for_stall_T_5 = 5'h2 == work_state ? _access_work_state_for_stall_T_1 : work_state; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_for_stall_T_7 = 5'h18 == work_state ? state_ready_lookup_should_be :
    _access_work_state_for_stall_T_5; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_for_stall_T_9 = 5'h5 == work_state ? _access_work_state_for_stall_T_3 :
    _access_work_state_for_stall_T_7; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_for_stall_T_11 = 5'h19 == work_state ? state_ready_lookup_should_be :
    _access_work_state_for_stall_T_9; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_for_stall_T_13 = 5'he == work_state ? 5'h18 : _access_work_state_for_stall_T_11; // @[Mux.scala 81:58]
  wire [4:0] access_work_state_for_stall = 5'h10 == work_state ? 5'h18 : _access_work_state_for_stall_T_13; // @[Mux.scala 81:58]
  wire  stage2_stall = access_work_state_for_stall[4:3] == 2'h3; // @[data_cache.scala 288:54]
  reg  stage2_sram_write_reg; // @[data_cache.scala 171:40]
  reg  stage1_stall_reg; // @[data_cache.scala 178:35]
  reg  write_access_complete_reg; // @[data_cache.scala 181:44]
  wire [2:0] _stage1_sram_size_reg_T_1 = io_sram_req ? io_sram_size : {{1'd0}, stage1_sram_size_reg}; // @[data_cache.scala 188:33]
  wire  _stage1_sram_req_reg_T_1 = stage2_stall ? 1'h0 : stage1_sram_req_reg; // @[data_cache.scala 190:60]
  wire [4:0] _state_lookup_for_less_delay_T_1 = 5'h18 == work_state ? state_ready_lookup_should_be : work_state; // @[Mux.scala 81:58]
  wire [4:0] state_lookup_for_less_delay = 5'h19 == work_state ? state_ready_lookup_should_be :
    _state_lookup_for_less_delay_T_1; // @[Mux.scala 81:58]
  wire  _way0_dirty_T = state_lookup_for_less_delay == 5'h19; // @[data_cache.scala 199:79]
  wire  _way0_dirty_T_2 = state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg; // @[data_cache.scala 199:96]
  wire  _way0_dirty_T_4 = state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
    stage1_sram_valid0_reg; // @[data_cache.scala 199:149]
  wire  _way0_dirty_T_5 = work_state == 5'he; // @[data_cache.scala 200:24]
  wire  _GEN_258 = 7'h1 == stage1_addr_line_mapping[10:4] ? lru_1 : lru_0; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_259 = 7'h2 == stage1_addr_line_mapping[10:4] ? lru_2 : _GEN_258; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_260 = 7'h3 == stage1_addr_line_mapping[10:4] ? lru_3 : _GEN_259; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_261 = 7'h4 == stage1_addr_line_mapping[10:4] ? lru_4 : _GEN_260; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_262 = 7'h5 == stage1_addr_line_mapping[10:4] ? lru_5 : _GEN_261; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_263 = 7'h6 == stage1_addr_line_mapping[10:4] ? lru_6 : _GEN_262; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_264 = 7'h7 == stage1_addr_line_mapping[10:4] ? lru_7 : _GEN_263; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_265 = 7'h8 == stage1_addr_line_mapping[10:4] ? lru_8 : _GEN_264; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_266 = 7'h9 == stage1_addr_line_mapping[10:4] ? lru_9 : _GEN_265; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_267 = 7'ha == stage1_addr_line_mapping[10:4] ? lru_10 : _GEN_266; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_268 = 7'hb == stage1_addr_line_mapping[10:4] ? lru_11 : _GEN_267; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_269 = 7'hc == stage1_addr_line_mapping[10:4] ? lru_12 : _GEN_268; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_270 = 7'hd == stage1_addr_line_mapping[10:4] ? lru_13 : _GEN_269; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_271 = 7'he == stage1_addr_line_mapping[10:4] ? lru_14 : _GEN_270; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_272 = 7'hf == stage1_addr_line_mapping[10:4] ? lru_15 : _GEN_271; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_273 = 7'h10 == stage1_addr_line_mapping[10:4] ? lru_16 : _GEN_272; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_274 = 7'h11 == stage1_addr_line_mapping[10:4] ? lru_17 : _GEN_273; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_275 = 7'h12 == stage1_addr_line_mapping[10:4] ? lru_18 : _GEN_274; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_276 = 7'h13 == stage1_addr_line_mapping[10:4] ? lru_19 : _GEN_275; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_277 = 7'h14 == stage1_addr_line_mapping[10:4] ? lru_20 : _GEN_276; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_278 = 7'h15 == stage1_addr_line_mapping[10:4] ? lru_21 : _GEN_277; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_279 = 7'h16 == stage1_addr_line_mapping[10:4] ? lru_22 : _GEN_278; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_280 = 7'h17 == stage1_addr_line_mapping[10:4] ? lru_23 : _GEN_279; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_281 = 7'h18 == stage1_addr_line_mapping[10:4] ? lru_24 : _GEN_280; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_282 = 7'h19 == stage1_addr_line_mapping[10:4] ? lru_25 : _GEN_281; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_283 = 7'h1a == stage1_addr_line_mapping[10:4] ? lru_26 : _GEN_282; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_284 = 7'h1b == stage1_addr_line_mapping[10:4] ? lru_27 : _GEN_283; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_285 = 7'h1c == stage1_addr_line_mapping[10:4] ? lru_28 : _GEN_284; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_286 = 7'h1d == stage1_addr_line_mapping[10:4] ? lru_29 : _GEN_285; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_287 = 7'h1e == stage1_addr_line_mapping[10:4] ? lru_30 : _GEN_286; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_288 = 7'h1f == stage1_addr_line_mapping[10:4] ? lru_31 : _GEN_287; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_289 = 7'h20 == stage1_addr_line_mapping[10:4] ? lru_32 : _GEN_288; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_290 = 7'h21 == stage1_addr_line_mapping[10:4] ? lru_33 : _GEN_289; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_291 = 7'h22 == stage1_addr_line_mapping[10:4] ? lru_34 : _GEN_290; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_292 = 7'h23 == stage1_addr_line_mapping[10:4] ? lru_35 : _GEN_291; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_293 = 7'h24 == stage1_addr_line_mapping[10:4] ? lru_36 : _GEN_292; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_294 = 7'h25 == stage1_addr_line_mapping[10:4] ? lru_37 : _GEN_293; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_295 = 7'h26 == stage1_addr_line_mapping[10:4] ? lru_38 : _GEN_294; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_296 = 7'h27 == stage1_addr_line_mapping[10:4] ? lru_39 : _GEN_295; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_297 = 7'h28 == stage1_addr_line_mapping[10:4] ? lru_40 : _GEN_296; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_298 = 7'h29 == stage1_addr_line_mapping[10:4] ? lru_41 : _GEN_297; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_299 = 7'h2a == stage1_addr_line_mapping[10:4] ? lru_42 : _GEN_298; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_300 = 7'h2b == stage1_addr_line_mapping[10:4] ? lru_43 : _GEN_299; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_301 = 7'h2c == stage1_addr_line_mapping[10:4] ? lru_44 : _GEN_300; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_302 = 7'h2d == stage1_addr_line_mapping[10:4] ? lru_45 : _GEN_301; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_303 = 7'h2e == stage1_addr_line_mapping[10:4] ? lru_46 : _GEN_302; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_304 = 7'h2f == stage1_addr_line_mapping[10:4] ? lru_47 : _GEN_303; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_305 = 7'h30 == stage1_addr_line_mapping[10:4] ? lru_48 : _GEN_304; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_306 = 7'h31 == stage1_addr_line_mapping[10:4] ? lru_49 : _GEN_305; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_307 = 7'h32 == stage1_addr_line_mapping[10:4] ? lru_50 : _GEN_306; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_308 = 7'h33 == stage1_addr_line_mapping[10:4] ? lru_51 : _GEN_307; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_309 = 7'h34 == stage1_addr_line_mapping[10:4] ? lru_52 : _GEN_308; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_310 = 7'h35 == stage1_addr_line_mapping[10:4] ? lru_53 : _GEN_309; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_311 = 7'h36 == stage1_addr_line_mapping[10:4] ? lru_54 : _GEN_310; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_312 = 7'h37 == stage1_addr_line_mapping[10:4] ? lru_55 : _GEN_311; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_313 = 7'h38 == stage1_addr_line_mapping[10:4] ? lru_56 : _GEN_312; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_314 = 7'h39 == stage1_addr_line_mapping[10:4] ? lru_57 : _GEN_313; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_315 = 7'h3a == stage1_addr_line_mapping[10:4] ? lru_58 : _GEN_314; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_316 = 7'h3b == stage1_addr_line_mapping[10:4] ? lru_59 : _GEN_315; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_317 = 7'h3c == stage1_addr_line_mapping[10:4] ? lru_60 : _GEN_316; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_318 = 7'h3d == stage1_addr_line_mapping[10:4] ? lru_61 : _GEN_317; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_319 = 7'h3e == stage1_addr_line_mapping[10:4] ? lru_62 : _GEN_318; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_320 = 7'h3f == stage1_addr_line_mapping[10:4] ? lru_63 : _GEN_319; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_321 = 7'h40 == stage1_addr_line_mapping[10:4] ? lru_64 : _GEN_320; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_322 = 7'h41 == stage1_addr_line_mapping[10:4] ? lru_65 : _GEN_321; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_323 = 7'h42 == stage1_addr_line_mapping[10:4] ? lru_66 : _GEN_322; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_324 = 7'h43 == stage1_addr_line_mapping[10:4] ? lru_67 : _GEN_323; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_325 = 7'h44 == stage1_addr_line_mapping[10:4] ? lru_68 : _GEN_324; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_326 = 7'h45 == stage1_addr_line_mapping[10:4] ? lru_69 : _GEN_325; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_327 = 7'h46 == stage1_addr_line_mapping[10:4] ? lru_70 : _GEN_326; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_328 = 7'h47 == stage1_addr_line_mapping[10:4] ? lru_71 : _GEN_327; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_329 = 7'h48 == stage1_addr_line_mapping[10:4] ? lru_72 : _GEN_328; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_330 = 7'h49 == stage1_addr_line_mapping[10:4] ? lru_73 : _GEN_329; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_331 = 7'h4a == stage1_addr_line_mapping[10:4] ? lru_74 : _GEN_330; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_332 = 7'h4b == stage1_addr_line_mapping[10:4] ? lru_75 : _GEN_331; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_333 = 7'h4c == stage1_addr_line_mapping[10:4] ? lru_76 : _GEN_332; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_334 = 7'h4d == stage1_addr_line_mapping[10:4] ? lru_77 : _GEN_333; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_335 = 7'h4e == stage1_addr_line_mapping[10:4] ? lru_78 : _GEN_334; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_336 = 7'h4f == stage1_addr_line_mapping[10:4] ? lru_79 : _GEN_335; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_337 = 7'h50 == stage1_addr_line_mapping[10:4] ? lru_80 : _GEN_336; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_338 = 7'h51 == stage1_addr_line_mapping[10:4] ? lru_81 : _GEN_337; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_339 = 7'h52 == stage1_addr_line_mapping[10:4] ? lru_82 : _GEN_338; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_340 = 7'h53 == stage1_addr_line_mapping[10:4] ? lru_83 : _GEN_339; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_341 = 7'h54 == stage1_addr_line_mapping[10:4] ? lru_84 : _GEN_340; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_342 = 7'h55 == stage1_addr_line_mapping[10:4] ? lru_85 : _GEN_341; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_343 = 7'h56 == stage1_addr_line_mapping[10:4] ? lru_86 : _GEN_342; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_344 = 7'h57 == stage1_addr_line_mapping[10:4] ? lru_87 : _GEN_343; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_345 = 7'h58 == stage1_addr_line_mapping[10:4] ? lru_88 : _GEN_344; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_346 = 7'h59 == stage1_addr_line_mapping[10:4] ? lru_89 : _GEN_345; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_347 = 7'h5a == stage1_addr_line_mapping[10:4] ? lru_90 : _GEN_346; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_348 = 7'h5b == stage1_addr_line_mapping[10:4] ? lru_91 : _GEN_347; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_349 = 7'h5c == stage1_addr_line_mapping[10:4] ? lru_92 : _GEN_348; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_350 = 7'h5d == stage1_addr_line_mapping[10:4] ? lru_93 : _GEN_349; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_351 = 7'h5e == stage1_addr_line_mapping[10:4] ? lru_94 : _GEN_350; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_352 = 7'h5f == stage1_addr_line_mapping[10:4] ? lru_95 : _GEN_351; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_353 = 7'h60 == stage1_addr_line_mapping[10:4] ? lru_96 : _GEN_352; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_354 = 7'h61 == stage1_addr_line_mapping[10:4] ? lru_97 : _GEN_353; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_355 = 7'h62 == stage1_addr_line_mapping[10:4] ? lru_98 : _GEN_354; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_356 = 7'h63 == stage1_addr_line_mapping[10:4] ? lru_99 : _GEN_355; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_357 = 7'h64 == stage1_addr_line_mapping[10:4] ? lru_100 : _GEN_356; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_358 = 7'h65 == stage1_addr_line_mapping[10:4] ? lru_101 : _GEN_357; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_359 = 7'h66 == stage1_addr_line_mapping[10:4] ? lru_102 : _GEN_358; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_360 = 7'h67 == stage1_addr_line_mapping[10:4] ? lru_103 : _GEN_359; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_361 = 7'h68 == stage1_addr_line_mapping[10:4] ? lru_104 : _GEN_360; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_362 = 7'h69 == stage1_addr_line_mapping[10:4] ? lru_105 : _GEN_361; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_363 = 7'h6a == stage1_addr_line_mapping[10:4] ? lru_106 : _GEN_362; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_364 = 7'h6b == stage1_addr_line_mapping[10:4] ? lru_107 : _GEN_363; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_365 = 7'h6c == stage1_addr_line_mapping[10:4] ? lru_108 : _GEN_364; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_366 = 7'h6d == stage1_addr_line_mapping[10:4] ? lru_109 : _GEN_365; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_367 = 7'h6e == stage1_addr_line_mapping[10:4] ? lru_110 : _GEN_366; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_368 = 7'h6f == stage1_addr_line_mapping[10:4] ? lru_111 : _GEN_367; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_369 = 7'h70 == stage1_addr_line_mapping[10:4] ? lru_112 : _GEN_368; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_370 = 7'h71 == stage1_addr_line_mapping[10:4] ? lru_113 : _GEN_369; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_371 = 7'h72 == stage1_addr_line_mapping[10:4] ? lru_114 : _GEN_370; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_372 = 7'h73 == stage1_addr_line_mapping[10:4] ? lru_115 : _GEN_371; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_373 = 7'h74 == stage1_addr_line_mapping[10:4] ? lru_116 : _GEN_372; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_374 = 7'h75 == stage1_addr_line_mapping[10:4] ? lru_117 : _GEN_373; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_375 = 7'h76 == stage1_addr_line_mapping[10:4] ? lru_118 : _GEN_374; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_376 = 7'h77 == stage1_addr_line_mapping[10:4] ? lru_119 : _GEN_375; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_377 = 7'h78 == stage1_addr_line_mapping[10:4] ? lru_120 : _GEN_376; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_378 = 7'h79 == stage1_addr_line_mapping[10:4] ? lru_121 : _GEN_377; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_379 = 7'h7a == stage1_addr_line_mapping[10:4] ? lru_122 : _GEN_378; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_380 = 7'h7b == stage1_addr_line_mapping[10:4] ? lru_123 : _GEN_379; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_381 = 7'h7c == stage1_addr_line_mapping[10:4] ? lru_124 : _GEN_380; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_382 = 7'h7d == stage1_addr_line_mapping[10:4] ? lru_125 : _GEN_381; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_383 = 7'h7e == stage1_addr_line_mapping[10:4] ? lru_126 : _GEN_382; // @[data_cache.scala 200:{86,86}]
  wire  _GEN_384 = 7'h7f == stage1_addr_line_mapping[10:4] ? lru_127 : _GEN_383; // @[data_cache.scala 200:{86,86}]
  wire  _way0_dirty_T_7 = ~_GEN_384; // @[data_cache.scala 200:86]
  wire  _way0_dirty_T_9 = work_state == 5'h10; // @[data_cache.scala 201:24]
  wire  _way0_dirty_T_12 = work_state == 5'h10 & _way0_dirty_T_7; // @[data_cache.scala 201:52]
  wire  _GEN_514 = 7'h1 == stage1_addr_line_mapping[10:4] ? way0_dirty_1 : way0_dirty_0; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_515 = 7'h2 == stage1_addr_line_mapping[10:4] ? way0_dirty_2 : _GEN_514; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_516 = 7'h3 == stage1_addr_line_mapping[10:4] ? way0_dirty_3 : _GEN_515; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_517 = 7'h4 == stage1_addr_line_mapping[10:4] ? way0_dirty_4 : _GEN_516; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_518 = 7'h5 == stage1_addr_line_mapping[10:4] ? way0_dirty_5 : _GEN_517; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_519 = 7'h6 == stage1_addr_line_mapping[10:4] ? way0_dirty_6 : _GEN_518; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_520 = 7'h7 == stage1_addr_line_mapping[10:4] ? way0_dirty_7 : _GEN_519; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_521 = 7'h8 == stage1_addr_line_mapping[10:4] ? way0_dirty_8 : _GEN_520; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_522 = 7'h9 == stage1_addr_line_mapping[10:4] ? way0_dirty_9 : _GEN_521; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_523 = 7'ha == stage1_addr_line_mapping[10:4] ? way0_dirty_10 : _GEN_522; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_524 = 7'hb == stage1_addr_line_mapping[10:4] ? way0_dirty_11 : _GEN_523; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_525 = 7'hc == stage1_addr_line_mapping[10:4] ? way0_dirty_12 : _GEN_524; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_526 = 7'hd == stage1_addr_line_mapping[10:4] ? way0_dirty_13 : _GEN_525; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_527 = 7'he == stage1_addr_line_mapping[10:4] ? way0_dirty_14 : _GEN_526; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_528 = 7'hf == stage1_addr_line_mapping[10:4] ? way0_dirty_15 : _GEN_527; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_529 = 7'h10 == stage1_addr_line_mapping[10:4] ? way0_dirty_16 : _GEN_528; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_530 = 7'h11 == stage1_addr_line_mapping[10:4] ? way0_dirty_17 : _GEN_529; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_531 = 7'h12 == stage1_addr_line_mapping[10:4] ? way0_dirty_18 : _GEN_530; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_532 = 7'h13 == stage1_addr_line_mapping[10:4] ? way0_dirty_19 : _GEN_531; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_533 = 7'h14 == stage1_addr_line_mapping[10:4] ? way0_dirty_20 : _GEN_532; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_534 = 7'h15 == stage1_addr_line_mapping[10:4] ? way0_dirty_21 : _GEN_533; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_535 = 7'h16 == stage1_addr_line_mapping[10:4] ? way0_dirty_22 : _GEN_534; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_536 = 7'h17 == stage1_addr_line_mapping[10:4] ? way0_dirty_23 : _GEN_535; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_537 = 7'h18 == stage1_addr_line_mapping[10:4] ? way0_dirty_24 : _GEN_536; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_538 = 7'h19 == stage1_addr_line_mapping[10:4] ? way0_dirty_25 : _GEN_537; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_539 = 7'h1a == stage1_addr_line_mapping[10:4] ? way0_dirty_26 : _GEN_538; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_540 = 7'h1b == stage1_addr_line_mapping[10:4] ? way0_dirty_27 : _GEN_539; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_541 = 7'h1c == stage1_addr_line_mapping[10:4] ? way0_dirty_28 : _GEN_540; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_542 = 7'h1d == stage1_addr_line_mapping[10:4] ? way0_dirty_29 : _GEN_541; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_543 = 7'h1e == stage1_addr_line_mapping[10:4] ? way0_dirty_30 : _GEN_542; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_544 = 7'h1f == stage1_addr_line_mapping[10:4] ? way0_dirty_31 : _GEN_543; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_545 = 7'h20 == stage1_addr_line_mapping[10:4] ? way0_dirty_32 : _GEN_544; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_546 = 7'h21 == stage1_addr_line_mapping[10:4] ? way0_dirty_33 : _GEN_545; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_547 = 7'h22 == stage1_addr_line_mapping[10:4] ? way0_dirty_34 : _GEN_546; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_548 = 7'h23 == stage1_addr_line_mapping[10:4] ? way0_dirty_35 : _GEN_547; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_549 = 7'h24 == stage1_addr_line_mapping[10:4] ? way0_dirty_36 : _GEN_548; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_550 = 7'h25 == stage1_addr_line_mapping[10:4] ? way0_dirty_37 : _GEN_549; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_551 = 7'h26 == stage1_addr_line_mapping[10:4] ? way0_dirty_38 : _GEN_550; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_552 = 7'h27 == stage1_addr_line_mapping[10:4] ? way0_dirty_39 : _GEN_551; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_553 = 7'h28 == stage1_addr_line_mapping[10:4] ? way0_dirty_40 : _GEN_552; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_554 = 7'h29 == stage1_addr_line_mapping[10:4] ? way0_dirty_41 : _GEN_553; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_555 = 7'h2a == stage1_addr_line_mapping[10:4] ? way0_dirty_42 : _GEN_554; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_556 = 7'h2b == stage1_addr_line_mapping[10:4] ? way0_dirty_43 : _GEN_555; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_557 = 7'h2c == stage1_addr_line_mapping[10:4] ? way0_dirty_44 : _GEN_556; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_558 = 7'h2d == stage1_addr_line_mapping[10:4] ? way0_dirty_45 : _GEN_557; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_559 = 7'h2e == stage1_addr_line_mapping[10:4] ? way0_dirty_46 : _GEN_558; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_560 = 7'h2f == stage1_addr_line_mapping[10:4] ? way0_dirty_47 : _GEN_559; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_561 = 7'h30 == stage1_addr_line_mapping[10:4] ? way0_dirty_48 : _GEN_560; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_562 = 7'h31 == stage1_addr_line_mapping[10:4] ? way0_dirty_49 : _GEN_561; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_563 = 7'h32 == stage1_addr_line_mapping[10:4] ? way0_dirty_50 : _GEN_562; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_564 = 7'h33 == stage1_addr_line_mapping[10:4] ? way0_dirty_51 : _GEN_563; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_565 = 7'h34 == stage1_addr_line_mapping[10:4] ? way0_dirty_52 : _GEN_564; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_566 = 7'h35 == stage1_addr_line_mapping[10:4] ? way0_dirty_53 : _GEN_565; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_567 = 7'h36 == stage1_addr_line_mapping[10:4] ? way0_dirty_54 : _GEN_566; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_568 = 7'h37 == stage1_addr_line_mapping[10:4] ? way0_dirty_55 : _GEN_567; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_569 = 7'h38 == stage1_addr_line_mapping[10:4] ? way0_dirty_56 : _GEN_568; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_570 = 7'h39 == stage1_addr_line_mapping[10:4] ? way0_dirty_57 : _GEN_569; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_571 = 7'h3a == stage1_addr_line_mapping[10:4] ? way0_dirty_58 : _GEN_570; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_572 = 7'h3b == stage1_addr_line_mapping[10:4] ? way0_dirty_59 : _GEN_571; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_573 = 7'h3c == stage1_addr_line_mapping[10:4] ? way0_dirty_60 : _GEN_572; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_574 = 7'h3d == stage1_addr_line_mapping[10:4] ? way0_dirty_61 : _GEN_573; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_575 = 7'h3e == stage1_addr_line_mapping[10:4] ? way0_dirty_62 : _GEN_574; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_576 = 7'h3f == stage1_addr_line_mapping[10:4] ? way0_dirty_63 : _GEN_575; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_577 = 7'h40 == stage1_addr_line_mapping[10:4] ? way0_dirty_64 : _GEN_576; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_578 = 7'h41 == stage1_addr_line_mapping[10:4] ? way0_dirty_65 : _GEN_577; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_579 = 7'h42 == stage1_addr_line_mapping[10:4] ? way0_dirty_66 : _GEN_578; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_580 = 7'h43 == stage1_addr_line_mapping[10:4] ? way0_dirty_67 : _GEN_579; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_581 = 7'h44 == stage1_addr_line_mapping[10:4] ? way0_dirty_68 : _GEN_580; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_582 = 7'h45 == stage1_addr_line_mapping[10:4] ? way0_dirty_69 : _GEN_581; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_583 = 7'h46 == stage1_addr_line_mapping[10:4] ? way0_dirty_70 : _GEN_582; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_584 = 7'h47 == stage1_addr_line_mapping[10:4] ? way0_dirty_71 : _GEN_583; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_585 = 7'h48 == stage1_addr_line_mapping[10:4] ? way0_dirty_72 : _GEN_584; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_586 = 7'h49 == stage1_addr_line_mapping[10:4] ? way0_dirty_73 : _GEN_585; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_587 = 7'h4a == stage1_addr_line_mapping[10:4] ? way0_dirty_74 : _GEN_586; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_588 = 7'h4b == stage1_addr_line_mapping[10:4] ? way0_dirty_75 : _GEN_587; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_589 = 7'h4c == stage1_addr_line_mapping[10:4] ? way0_dirty_76 : _GEN_588; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_590 = 7'h4d == stage1_addr_line_mapping[10:4] ? way0_dirty_77 : _GEN_589; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_591 = 7'h4e == stage1_addr_line_mapping[10:4] ? way0_dirty_78 : _GEN_590; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_592 = 7'h4f == stage1_addr_line_mapping[10:4] ? way0_dirty_79 : _GEN_591; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_593 = 7'h50 == stage1_addr_line_mapping[10:4] ? way0_dirty_80 : _GEN_592; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_594 = 7'h51 == stage1_addr_line_mapping[10:4] ? way0_dirty_81 : _GEN_593; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_595 = 7'h52 == stage1_addr_line_mapping[10:4] ? way0_dirty_82 : _GEN_594; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_596 = 7'h53 == stage1_addr_line_mapping[10:4] ? way0_dirty_83 : _GEN_595; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_597 = 7'h54 == stage1_addr_line_mapping[10:4] ? way0_dirty_84 : _GEN_596; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_598 = 7'h55 == stage1_addr_line_mapping[10:4] ? way0_dirty_85 : _GEN_597; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_599 = 7'h56 == stage1_addr_line_mapping[10:4] ? way0_dirty_86 : _GEN_598; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_600 = 7'h57 == stage1_addr_line_mapping[10:4] ? way0_dirty_87 : _GEN_599; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_601 = 7'h58 == stage1_addr_line_mapping[10:4] ? way0_dirty_88 : _GEN_600; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_602 = 7'h59 == stage1_addr_line_mapping[10:4] ? way0_dirty_89 : _GEN_601; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_603 = 7'h5a == stage1_addr_line_mapping[10:4] ? way0_dirty_90 : _GEN_602; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_604 = 7'h5b == stage1_addr_line_mapping[10:4] ? way0_dirty_91 : _GEN_603; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_605 = 7'h5c == stage1_addr_line_mapping[10:4] ? way0_dirty_92 : _GEN_604; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_606 = 7'h5d == stage1_addr_line_mapping[10:4] ? way0_dirty_93 : _GEN_605; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_607 = 7'h5e == stage1_addr_line_mapping[10:4] ? way0_dirty_94 : _GEN_606; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_608 = 7'h5f == stage1_addr_line_mapping[10:4] ? way0_dirty_95 : _GEN_607; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_609 = 7'h60 == stage1_addr_line_mapping[10:4] ? way0_dirty_96 : _GEN_608; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_610 = 7'h61 == stage1_addr_line_mapping[10:4] ? way0_dirty_97 : _GEN_609; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_611 = 7'h62 == stage1_addr_line_mapping[10:4] ? way0_dirty_98 : _GEN_610; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_612 = 7'h63 == stage1_addr_line_mapping[10:4] ? way0_dirty_99 : _GEN_611; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_613 = 7'h64 == stage1_addr_line_mapping[10:4] ? way0_dirty_100 : _GEN_612; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_614 = 7'h65 == stage1_addr_line_mapping[10:4] ? way0_dirty_101 : _GEN_613; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_615 = 7'h66 == stage1_addr_line_mapping[10:4] ? way0_dirty_102 : _GEN_614; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_616 = 7'h67 == stage1_addr_line_mapping[10:4] ? way0_dirty_103 : _GEN_615; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_617 = 7'h68 == stage1_addr_line_mapping[10:4] ? way0_dirty_104 : _GEN_616; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_618 = 7'h69 == stage1_addr_line_mapping[10:4] ? way0_dirty_105 : _GEN_617; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_619 = 7'h6a == stage1_addr_line_mapping[10:4] ? way0_dirty_106 : _GEN_618; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_620 = 7'h6b == stage1_addr_line_mapping[10:4] ? way0_dirty_107 : _GEN_619; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_621 = 7'h6c == stage1_addr_line_mapping[10:4] ? way0_dirty_108 : _GEN_620; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_622 = 7'h6d == stage1_addr_line_mapping[10:4] ? way0_dirty_109 : _GEN_621; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_623 = 7'h6e == stage1_addr_line_mapping[10:4] ? way0_dirty_110 : _GEN_622; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_624 = 7'h6f == stage1_addr_line_mapping[10:4] ? way0_dirty_111 : _GEN_623; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_625 = 7'h70 == stage1_addr_line_mapping[10:4] ? way0_dirty_112 : _GEN_624; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_626 = 7'h71 == stage1_addr_line_mapping[10:4] ? way0_dirty_113 : _GEN_625; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_627 = 7'h72 == stage1_addr_line_mapping[10:4] ? way0_dirty_114 : _GEN_626; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_628 = 7'h73 == stage1_addr_line_mapping[10:4] ? way0_dirty_115 : _GEN_627; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_629 = 7'h74 == stage1_addr_line_mapping[10:4] ? way0_dirty_116 : _GEN_628; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_630 = 7'h75 == stage1_addr_line_mapping[10:4] ? way0_dirty_117 : _GEN_629; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_631 = 7'h76 == stage1_addr_line_mapping[10:4] ? way0_dirty_118 : _GEN_630; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_632 = 7'h77 == stage1_addr_line_mapping[10:4] ? way0_dirty_119 : _GEN_631; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_633 = 7'h78 == stage1_addr_line_mapping[10:4] ? way0_dirty_120 : _GEN_632; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_634 = 7'h79 == stage1_addr_line_mapping[10:4] ? way0_dirty_121 : _GEN_633; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_635 = 7'h7a == stage1_addr_line_mapping[10:4] ? way0_dirty_122 : _GEN_634; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_636 = 7'h7b == stage1_addr_line_mapping[10:4] ? way0_dirty_123 : _GEN_635; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_637 = 7'h7c == stage1_addr_line_mapping[10:4] ? way0_dirty_124 : _GEN_636; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_638 = 7'h7d == stage1_addr_line_mapping[10:4] ? way0_dirty_125 : _GEN_637; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_639 = 7'h7e == stage1_addr_line_mapping[10:4] ? way0_dirty_126 : _GEN_638; // @[data_cache.scala 201:{12,12}]
  wire  _GEN_640 = 7'h7f == stage1_addr_line_mapping[10:4] ? way0_dirty_127 : _GEN_639; // @[data_cache.scala 201:{12,12}]
  wire  _way0_dirty_T_14 = work_state == 5'h10 & _way0_dirty_T_7 | _GEN_640; // @[data_cache.scala 201:12]
  wire  _way0_dirty_T_15 = work_state == 5'he & ~_GEN_384 ? 1'h0 : _way0_dirty_T_14; // @[data_cache.scala 200:12]
  wire  _way1_dirty_T_4 = _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg; // @[data_cache.scala 203:149]
  wire  _way1_dirty_T_12 = _way0_dirty_T_9 & _GEN_384; // @[data_cache.scala 205:52]
  wire  _GEN_1026 = 7'h1 == stage1_addr_line_mapping[10:4] ? way1_dirty_1 : way1_dirty_0; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1027 = 7'h2 == stage1_addr_line_mapping[10:4] ? way1_dirty_2 : _GEN_1026; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1028 = 7'h3 == stage1_addr_line_mapping[10:4] ? way1_dirty_3 : _GEN_1027; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1029 = 7'h4 == stage1_addr_line_mapping[10:4] ? way1_dirty_4 : _GEN_1028; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1030 = 7'h5 == stage1_addr_line_mapping[10:4] ? way1_dirty_5 : _GEN_1029; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1031 = 7'h6 == stage1_addr_line_mapping[10:4] ? way1_dirty_6 : _GEN_1030; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1032 = 7'h7 == stage1_addr_line_mapping[10:4] ? way1_dirty_7 : _GEN_1031; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1033 = 7'h8 == stage1_addr_line_mapping[10:4] ? way1_dirty_8 : _GEN_1032; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1034 = 7'h9 == stage1_addr_line_mapping[10:4] ? way1_dirty_9 : _GEN_1033; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1035 = 7'ha == stage1_addr_line_mapping[10:4] ? way1_dirty_10 : _GEN_1034; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1036 = 7'hb == stage1_addr_line_mapping[10:4] ? way1_dirty_11 : _GEN_1035; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1037 = 7'hc == stage1_addr_line_mapping[10:4] ? way1_dirty_12 : _GEN_1036; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1038 = 7'hd == stage1_addr_line_mapping[10:4] ? way1_dirty_13 : _GEN_1037; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1039 = 7'he == stage1_addr_line_mapping[10:4] ? way1_dirty_14 : _GEN_1038; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1040 = 7'hf == stage1_addr_line_mapping[10:4] ? way1_dirty_15 : _GEN_1039; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1041 = 7'h10 == stage1_addr_line_mapping[10:4] ? way1_dirty_16 : _GEN_1040; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1042 = 7'h11 == stage1_addr_line_mapping[10:4] ? way1_dirty_17 : _GEN_1041; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1043 = 7'h12 == stage1_addr_line_mapping[10:4] ? way1_dirty_18 : _GEN_1042; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1044 = 7'h13 == stage1_addr_line_mapping[10:4] ? way1_dirty_19 : _GEN_1043; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1045 = 7'h14 == stage1_addr_line_mapping[10:4] ? way1_dirty_20 : _GEN_1044; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1046 = 7'h15 == stage1_addr_line_mapping[10:4] ? way1_dirty_21 : _GEN_1045; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1047 = 7'h16 == stage1_addr_line_mapping[10:4] ? way1_dirty_22 : _GEN_1046; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1048 = 7'h17 == stage1_addr_line_mapping[10:4] ? way1_dirty_23 : _GEN_1047; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1049 = 7'h18 == stage1_addr_line_mapping[10:4] ? way1_dirty_24 : _GEN_1048; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1050 = 7'h19 == stage1_addr_line_mapping[10:4] ? way1_dirty_25 : _GEN_1049; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1051 = 7'h1a == stage1_addr_line_mapping[10:4] ? way1_dirty_26 : _GEN_1050; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1052 = 7'h1b == stage1_addr_line_mapping[10:4] ? way1_dirty_27 : _GEN_1051; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1053 = 7'h1c == stage1_addr_line_mapping[10:4] ? way1_dirty_28 : _GEN_1052; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1054 = 7'h1d == stage1_addr_line_mapping[10:4] ? way1_dirty_29 : _GEN_1053; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1055 = 7'h1e == stage1_addr_line_mapping[10:4] ? way1_dirty_30 : _GEN_1054; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1056 = 7'h1f == stage1_addr_line_mapping[10:4] ? way1_dirty_31 : _GEN_1055; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1057 = 7'h20 == stage1_addr_line_mapping[10:4] ? way1_dirty_32 : _GEN_1056; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1058 = 7'h21 == stage1_addr_line_mapping[10:4] ? way1_dirty_33 : _GEN_1057; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1059 = 7'h22 == stage1_addr_line_mapping[10:4] ? way1_dirty_34 : _GEN_1058; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1060 = 7'h23 == stage1_addr_line_mapping[10:4] ? way1_dirty_35 : _GEN_1059; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1061 = 7'h24 == stage1_addr_line_mapping[10:4] ? way1_dirty_36 : _GEN_1060; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1062 = 7'h25 == stage1_addr_line_mapping[10:4] ? way1_dirty_37 : _GEN_1061; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1063 = 7'h26 == stage1_addr_line_mapping[10:4] ? way1_dirty_38 : _GEN_1062; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1064 = 7'h27 == stage1_addr_line_mapping[10:4] ? way1_dirty_39 : _GEN_1063; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1065 = 7'h28 == stage1_addr_line_mapping[10:4] ? way1_dirty_40 : _GEN_1064; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1066 = 7'h29 == stage1_addr_line_mapping[10:4] ? way1_dirty_41 : _GEN_1065; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1067 = 7'h2a == stage1_addr_line_mapping[10:4] ? way1_dirty_42 : _GEN_1066; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1068 = 7'h2b == stage1_addr_line_mapping[10:4] ? way1_dirty_43 : _GEN_1067; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1069 = 7'h2c == stage1_addr_line_mapping[10:4] ? way1_dirty_44 : _GEN_1068; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1070 = 7'h2d == stage1_addr_line_mapping[10:4] ? way1_dirty_45 : _GEN_1069; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1071 = 7'h2e == stage1_addr_line_mapping[10:4] ? way1_dirty_46 : _GEN_1070; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1072 = 7'h2f == stage1_addr_line_mapping[10:4] ? way1_dirty_47 : _GEN_1071; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1073 = 7'h30 == stage1_addr_line_mapping[10:4] ? way1_dirty_48 : _GEN_1072; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1074 = 7'h31 == stage1_addr_line_mapping[10:4] ? way1_dirty_49 : _GEN_1073; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1075 = 7'h32 == stage1_addr_line_mapping[10:4] ? way1_dirty_50 : _GEN_1074; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1076 = 7'h33 == stage1_addr_line_mapping[10:4] ? way1_dirty_51 : _GEN_1075; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1077 = 7'h34 == stage1_addr_line_mapping[10:4] ? way1_dirty_52 : _GEN_1076; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1078 = 7'h35 == stage1_addr_line_mapping[10:4] ? way1_dirty_53 : _GEN_1077; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1079 = 7'h36 == stage1_addr_line_mapping[10:4] ? way1_dirty_54 : _GEN_1078; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1080 = 7'h37 == stage1_addr_line_mapping[10:4] ? way1_dirty_55 : _GEN_1079; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1081 = 7'h38 == stage1_addr_line_mapping[10:4] ? way1_dirty_56 : _GEN_1080; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1082 = 7'h39 == stage1_addr_line_mapping[10:4] ? way1_dirty_57 : _GEN_1081; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1083 = 7'h3a == stage1_addr_line_mapping[10:4] ? way1_dirty_58 : _GEN_1082; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1084 = 7'h3b == stage1_addr_line_mapping[10:4] ? way1_dirty_59 : _GEN_1083; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1085 = 7'h3c == stage1_addr_line_mapping[10:4] ? way1_dirty_60 : _GEN_1084; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1086 = 7'h3d == stage1_addr_line_mapping[10:4] ? way1_dirty_61 : _GEN_1085; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1087 = 7'h3e == stage1_addr_line_mapping[10:4] ? way1_dirty_62 : _GEN_1086; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1088 = 7'h3f == stage1_addr_line_mapping[10:4] ? way1_dirty_63 : _GEN_1087; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1089 = 7'h40 == stage1_addr_line_mapping[10:4] ? way1_dirty_64 : _GEN_1088; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1090 = 7'h41 == stage1_addr_line_mapping[10:4] ? way1_dirty_65 : _GEN_1089; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1091 = 7'h42 == stage1_addr_line_mapping[10:4] ? way1_dirty_66 : _GEN_1090; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1092 = 7'h43 == stage1_addr_line_mapping[10:4] ? way1_dirty_67 : _GEN_1091; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1093 = 7'h44 == stage1_addr_line_mapping[10:4] ? way1_dirty_68 : _GEN_1092; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1094 = 7'h45 == stage1_addr_line_mapping[10:4] ? way1_dirty_69 : _GEN_1093; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1095 = 7'h46 == stage1_addr_line_mapping[10:4] ? way1_dirty_70 : _GEN_1094; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1096 = 7'h47 == stage1_addr_line_mapping[10:4] ? way1_dirty_71 : _GEN_1095; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1097 = 7'h48 == stage1_addr_line_mapping[10:4] ? way1_dirty_72 : _GEN_1096; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1098 = 7'h49 == stage1_addr_line_mapping[10:4] ? way1_dirty_73 : _GEN_1097; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1099 = 7'h4a == stage1_addr_line_mapping[10:4] ? way1_dirty_74 : _GEN_1098; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1100 = 7'h4b == stage1_addr_line_mapping[10:4] ? way1_dirty_75 : _GEN_1099; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1101 = 7'h4c == stage1_addr_line_mapping[10:4] ? way1_dirty_76 : _GEN_1100; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1102 = 7'h4d == stage1_addr_line_mapping[10:4] ? way1_dirty_77 : _GEN_1101; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1103 = 7'h4e == stage1_addr_line_mapping[10:4] ? way1_dirty_78 : _GEN_1102; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1104 = 7'h4f == stage1_addr_line_mapping[10:4] ? way1_dirty_79 : _GEN_1103; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1105 = 7'h50 == stage1_addr_line_mapping[10:4] ? way1_dirty_80 : _GEN_1104; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1106 = 7'h51 == stage1_addr_line_mapping[10:4] ? way1_dirty_81 : _GEN_1105; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1107 = 7'h52 == stage1_addr_line_mapping[10:4] ? way1_dirty_82 : _GEN_1106; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1108 = 7'h53 == stage1_addr_line_mapping[10:4] ? way1_dirty_83 : _GEN_1107; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1109 = 7'h54 == stage1_addr_line_mapping[10:4] ? way1_dirty_84 : _GEN_1108; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1110 = 7'h55 == stage1_addr_line_mapping[10:4] ? way1_dirty_85 : _GEN_1109; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1111 = 7'h56 == stage1_addr_line_mapping[10:4] ? way1_dirty_86 : _GEN_1110; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1112 = 7'h57 == stage1_addr_line_mapping[10:4] ? way1_dirty_87 : _GEN_1111; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1113 = 7'h58 == stage1_addr_line_mapping[10:4] ? way1_dirty_88 : _GEN_1112; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1114 = 7'h59 == stage1_addr_line_mapping[10:4] ? way1_dirty_89 : _GEN_1113; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1115 = 7'h5a == stage1_addr_line_mapping[10:4] ? way1_dirty_90 : _GEN_1114; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1116 = 7'h5b == stage1_addr_line_mapping[10:4] ? way1_dirty_91 : _GEN_1115; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1117 = 7'h5c == stage1_addr_line_mapping[10:4] ? way1_dirty_92 : _GEN_1116; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1118 = 7'h5d == stage1_addr_line_mapping[10:4] ? way1_dirty_93 : _GEN_1117; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1119 = 7'h5e == stage1_addr_line_mapping[10:4] ? way1_dirty_94 : _GEN_1118; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1120 = 7'h5f == stage1_addr_line_mapping[10:4] ? way1_dirty_95 : _GEN_1119; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1121 = 7'h60 == stage1_addr_line_mapping[10:4] ? way1_dirty_96 : _GEN_1120; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1122 = 7'h61 == stage1_addr_line_mapping[10:4] ? way1_dirty_97 : _GEN_1121; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1123 = 7'h62 == stage1_addr_line_mapping[10:4] ? way1_dirty_98 : _GEN_1122; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1124 = 7'h63 == stage1_addr_line_mapping[10:4] ? way1_dirty_99 : _GEN_1123; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1125 = 7'h64 == stage1_addr_line_mapping[10:4] ? way1_dirty_100 : _GEN_1124; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1126 = 7'h65 == stage1_addr_line_mapping[10:4] ? way1_dirty_101 : _GEN_1125; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1127 = 7'h66 == stage1_addr_line_mapping[10:4] ? way1_dirty_102 : _GEN_1126; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1128 = 7'h67 == stage1_addr_line_mapping[10:4] ? way1_dirty_103 : _GEN_1127; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1129 = 7'h68 == stage1_addr_line_mapping[10:4] ? way1_dirty_104 : _GEN_1128; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1130 = 7'h69 == stage1_addr_line_mapping[10:4] ? way1_dirty_105 : _GEN_1129; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1131 = 7'h6a == stage1_addr_line_mapping[10:4] ? way1_dirty_106 : _GEN_1130; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1132 = 7'h6b == stage1_addr_line_mapping[10:4] ? way1_dirty_107 : _GEN_1131; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1133 = 7'h6c == stage1_addr_line_mapping[10:4] ? way1_dirty_108 : _GEN_1132; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1134 = 7'h6d == stage1_addr_line_mapping[10:4] ? way1_dirty_109 : _GEN_1133; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1135 = 7'h6e == stage1_addr_line_mapping[10:4] ? way1_dirty_110 : _GEN_1134; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1136 = 7'h6f == stage1_addr_line_mapping[10:4] ? way1_dirty_111 : _GEN_1135; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1137 = 7'h70 == stage1_addr_line_mapping[10:4] ? way1_dirty_112 : _GEN_1136; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1138 = 7'h71 == stage1_addr_line_mapping[10:4] ? way1_dirty_113 : _GEN_1137; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1139 = 7'h72 == stage1_addr_line_mapping[10:4] ? way1_dirty_114 : _GEN_1138; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1140 = 7'h73 == stage1_addr_line_mapping[10:4] ? way1_dirty_115 : _GEN_1139; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1141 = 7'h74 == stage1_addr_line_mapping[10:4] ? way1_dirty_116 : _GEN_1140; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1142 = 7'h75 == stage1_addr_line_mapping[10:4] ? way1_dirty_117 : _GEN_1141; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1143 = 7'h76 == stage1_addr_line_mapping[10:4] ? way1_dirty_118 : _GEN_1142; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1144 = 7'h77 == stage1_addr_line_mapping[10:4] ? way1_dirty_119 : _GEN_1143; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1145 = 7'h78 == stage1_addr_line_mapping[10:4] ? way1_dirty_120 : _GEN_1144; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1146 = 7'h79 == stage1_addr_line_mapping[10:4] ? way1_dirty_121 : _GEN_1145; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1147 = 7'h7a == stage1_addr_line_mapping[10:4] ? way1_dirty_122 : _GEN_1146; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1148 = 7'h7b == stage1_addr_line_mapping[10:4] ? way1_dirty_123 : _GEN_1147; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1149 = 7'h7c == stage1_addr_line_mapping[10:4] ? way1_dirty_124 : _GEN_1148; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1150 = 7'h7d == stage1_addr_line_mapping[10:4] ? way1_dirty_125 : _GEN_1149; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1151 = 7'h7e == stage1_addr_line_mapping[10:4] ? way1_dirty_126 : _GEN_1150; // @[data_cache.scala 205:{12,12}]
  wire  _GEN_1152 = 7'h7f == stage1_addr_line_mapping[10:4] ? way1_dirty_127 : _GEN_1151; // @[data_cache.scala 205:{12,12}]
  wire  _way1_dirty_T_14 = _way0_dirty_T_9 & _GEN_384 | _GEN_1152; // @[data_cache.scala 205:12]
  wire  _way1_dirty_T_15 = _way0_dirty_T_5 & _GEN_384 ? 1'h0 : _way1_dirty_T_14; // @[data_cache.scala 204:12]
  wire  dirty_victim = _way0_dirty_T_7 ? _GEN_640 : _GEN_1152; // @[data_cache.scala 209:24]
  wire [10:0] _T_3 = {data_write_back_counter[6:0],4'h0}; // @[Cat.scala 31:58]
  wire  _io_tlb_req_T_4 = ~stage1_addr_line_mapping[31] | stage1_addr_line_mapping[31:30] == 2'h3; // @[macros.scala 484:18]
  wire  _lru_T_4 = _hit_T_1 ? 1'h0 : _GEN_384; // @[data_cache.scala 230:12]
  wire  _lru_T_5 = _hit_T | _lru_T_4; // @[data_cache.scala 229:12]
  wire  _data_cache_under_write_all_back_T = work_state == 5'h18; // @[data_cache.scala 237:55]
  wire  _data_cache_under_write_all_back_T_1 = work_state == 5'h19; // @[data_cache.scala 237:90]
  wire [4:0] _state_ready_lookup_will_to_be_T_3 = stage1_sram_cache_reg ? 5'h19 : 5'h3; // @[data_cache.scala 240:16]
  wire [4:0] _state_ready_lookup_will_to_be_T_5 = stage1_sram_cache_reg ? 5'h19 : 5'h1; // @[data_cache.scala 240:88]
  wire [4:0] _state_ready_lookup_will_to_be_T_6 = stage1_sram_wr_reg ? _state_ready_lookup_will_to_be_T_3 :
    _state_ready_lookup_will_to_be_T_5; // @[data_cache.scala 239:55]
  wire [4:0] _state_ready_lookup_will_to_be_T_7 = stage1_sram_req_reg ? _state_ready_lookup_will_to_be_T_6 : 5'h19; // @[data_cache.scala 239:24]
  wire [1:0] _state_ready_lookup_will_to_be_T_12 = stage1_sram_wr_reg ? 2'h3 : 2'h1; // @[data_cache.scala 241:81]
  wire [3:0] _state_ready_lookup_will_to_be_T_15 = stage1_sram_wr_reg ? 4'h8 : 4'hc; // @[data_cache.scala 242:64]
  wire [3:0] _state_ready_lookup_will_to_be_T_16 = dirty_victim ? 4'h9 : _state_ready_lookup_will_to_be_T_15; // @[data_cache.scala 242:16]
  wire [3:0] _state_ready_lookup_will_to_be_T_17 = ~stage1_sram_cache_reg ? {{2'd0}, _state_ready_lookup_will_to_be_T_12
    } : _state_ready_lookup_will_to_be_T_16; // @[data_cache.scala 241:47]
  wire [4:0] _state_ready_lookup_will_to_be_T_18 = stage1_sram_req_reg ? {{1'd0}, _state_ready_lookup_will_to_be_T_17}
     : 5'h19; // @[data_cache.scala 241:16]
  wire [4:0] _state_ready_lookup_will_to_be_T_19 = hit ? _state_ready_lookup_will_to_be_T_7 :
    _state_ready_lookup_will_to_be_T_18; // @[data_cache.scala 239:16]
  wire [4:0] state_ready_lookup_will_to_be = io_fence_i_control ? 5'h11 : _state_ready_lookup_will_to_be_T_19; // @[data_cache.scala 238:41]
  wire [4:0] _access_work_state_T_1 = io_port_arready ? 5'h2 : work_state; // @[data_cache.scala 249:39]
  wire [2:0] _access_work_state_T_6 = io_port_wready ? 3'h5 : 3'h4; // @[data_cache.scala 252:66]
  wire [4:0] _access_work_state_T_7 = io_port_awready ? {{2'd0}, _access_work_state_T_6} : work_state; // @[data_cache.scala 252:39]
  wire [4:0] _access_work_state_T_9 = io_port_wready ? 5'h5 : work_state; // @[data_cache.scala 253:39]
  wire [4:0] _access_work_state_T_13 = io_port_arready ? 5'hd : work_state; // @[data_cache.scala 256:44]
  wire [4:0] _access_work_state_T_18 = stage1_sram_wr_reg ? 5'h10 : 5'he; // @[data_cache.scala 257:94]
  wire [4:0] _access_work_state_T_19 = io_port_rlast & io_port_rvalid ? _access_work_state_T_18 : work_state; // @[data_cache.scala 257:44]
  wire [4:0] _access_work_state_T_21 = io_port_awready ? 5'ha : work_state; // @[data_cache.scala 259:41]
  wire  _access_work_state_T_23 = write_counter == 3'h1; // @[data_cache.scala 260:81]
  wire  _access_work_state_T_24 = io_port_wready & write_counter == 3'h1; // @[data_cache.scala 260:64]
  wire [4:0] _access_work_state_T_25 = io_port_wready & write_counter == 3'h1 ? 5'hb : work_state; // @[data_cache.scala 260:41]
  wire [4:0] _access_work_state_T_27 = io_port_bvalid ? 5'hc : work_state; // @[data_cache.scala 261:41]
  wire [4:0] _access_work_state_T_29 = io_port_arready ? 5'h0 : work_state; // @[data_cache.scala 263:44]
  wire  _access_work_state_T_32 = io_port_rvalid & io_port_rlast; // @[data_cache.scala 264:68]
  wire [4:0] _access_work_state_T_33 = io_port_rvalid & io_port_rlast ? 5'h10 : work_state; // @[data_cache.scala 264:44]
  wire [4:0] _access_work_state_T_35 = io_port_awready ? 5'h6 : work_state; // @[data_cache.scala 266:41]
  wire [4:0] _access_work_state_T_39 = _access_work_state_T_24 ? 5'h7 : work_state; // @[data_cache.scala 267:41]
  wire [4:0] _access_work_state_T_41 = io_port_bvalid ? 5'h8 : work_state; // @[data_cache.scala 268:41]
  wire [4:0] _access_work_state_T_42 = data_all_write_back ? 5'h15 : work_state; // @[data_cache.scala 270:94]
  wire [4:0] _access_work_state_T_43 = data_should_write_back ? 5'h12 : _access_work_state_T_42; // @[data_cache.scala 270:41]
  wire [4:0] _access_work_state_T_45 = io_port_awready ? 5'h13 : work_state; // @[data_cache.scala 271:41]
  wire [4:0] _access_work_state_T_54 = 5'h1 == work_state ? _access_work_state_T_1 : work_state; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_56 = 5'h2 == work_state ? _access_work_state_for_stall_T_1 : _access_work_state_T_54; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_58 = 5'h18 == work_state ? state_ready_lookup_will_to_be : _access_work_state_T_56; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_60 = 5'h3 == work_state ? _access_work_state_T_7 : _access_work_state_T_58; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_62 = 5'h4 == work_state ? _access_work_state_T_9 : _access_work_state_T_60; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_64 = 5'h5 == work_state ? _access_work_state_for_stall_T_3 : _access_work_state_T_62; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_66 = 5'h19 == work_state ? state_ready_lookup_will_to_be : _access_work_state_T_64; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_68 = 5'hc == work_state ? _access_work_state_T_13 : _access_work_state_T_66; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_70 = 5'hd == work_state ? _access_work_state_T_19 : _access_work_state_T_68; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_72 = 5'he == work_state ? 5'h18 : _access_work_state_T_70; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_74 = 5'h9 == work_state ? _access_work_state_T_21 : _access_work_state_T_72; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_76 = 5'ha == work_state ? _access_work_state_T_25 : _access_work_state_T_74; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_78 = 5'hb == work_state ? _access_work_state_T_27 : _access_work_state_T_76; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_80 = 5'h8 == work_state ? _access_work_state_T_29 : _access_work_state_T_78; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_82 = 5'h0 == work_state ? _access_work_state_T_33 : _access_work_state_T_80; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_84 = 5'h10 == work_state ? 5'h18 : _access_work_state_T_82; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_86 = 5'hf == work_state ? _access_work_state_T_35 : _access_work_state_T_84; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_88 = 5'h6 == work_state ? _access_work_state_T_39 : _access_work_state_T_86; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_90 = 5'h7 == work_state ? _access_work_state_T_41 : _access_work_state_T_88; // @[Mux.scala 81:58]
  wire [4:0] _access_work_state_T_92 = 5'h11 == work_state ? _access_work_state_T_43 : _access_work_state_T_90; // @[Mux.scala 81:58]
  wire  _wait_data_T_3 = work_state == 5'hd; // @[data_cache.scala 293:24]
  wire [2:0] _GEN_3468 = {{2'd0}, stage1_addr_line_mapping[3]}; // @[data_cache.scala 293:98]
  wire  _write_counter_T = work_state == 5'ha; // @[data_cache.scala 295:37]
  wire  _write_counter_T_1 = work_state == 5'h9; // @[data_cache.scala 295:79]
  wire  _write_counter_T_2 = work_state == 5'ha | work_state == 5'h9; // @[data_cache.scala 295:65]
  wire [2:0] _write_counter_T_6 = write_counter + 3'h1; // @[data_cache.scala 295:190]
  wire [2:0] _write_counter_T_7 = _access_work_state_T_23 ? 3'h0 : _write_counter_T_6; // @[data_cache.scala 295:137]
  wire [2:0] _write_counter_T_8 = io_port_wready ? _write_counter_T_7 : write_counter; // @[data_cache.scala 295:111]
  wire  _write_counter_T_9 = work_state == 5'h6; // @[data_cache.scala 296:24]
  wire  _write_counter_T_10 = work_state == 5'hf; // @[data_cache.scala 296:67]
  wire [2:0] _read_counter_T_6 = read_counter + 3'h1; // @[data_cache.scala 298:163]
  wire [2:0] _read_counter_T_7 = io_port_rvalid ? _read_counter_T_6 : read_counter; // @[data_cache.scala 298:128]
  wire [2:0] _read_counter_T_8 = _access_work_state_T_32 ? 3'h0 : _read_counter_T_7; // @[data_cache.scala 298:72]
  wire  _read_counter_T_9 = work_state == 5'h0; // @[data_cache.scala 299:24]
  reg [63:0] stage2_sram_addr_reg; // @[Reg.scala 28:20]
  reg  stage2_hit0_reg; // @[data_cache.scala 321:34]
  wire [63:0] dcache_data_way0_0_rdata = dcache_data_io_rdata; // @[data_cache.scala 93:{36,36}]
  wire [63:0] dcache_data_way0_1_rdata = dcache_data_1_io_rdata; // @[data_cache.scala 93:{36,36}]
  wire [63:0] _GEN_2179 = stage2_sram_addr_reg[3] ? dcache_data_way0_1_rdata : dcache_data_way0_0_rdata; // @[data_cache.scala 346:{23,23}]
  wire [63:0] dcache_data_way1_0_rdata = dcache_data_2_io_rdata; // @[data_cache.scala 94:{36,36}]
  wire [63:0] dcache_data_way1_1_rdata = dcache_data_3_io_rdata; // @[data_cache.scala 94:{36,36}]
  wire [63:0] _GEN_2181 = stage2_sram_addr_reg[3] ? dcache_data_way1_1_rdata : dcache_data_way1_0_rdata; // @[data_cache.scala 346:{23,23}]
  wire [63:0] hit_word = stage2_hit0_reg ? _GEN_2179 : _GEN_2181; // @[data_cache.scala 346:23]
  wire [63:0] _GEN_2183 = write_counter[0] ? dcache_data_way1_1_rdata : dcache_data_way1_0_rdata; // @[data_cache.scala 356:{29,29}]
  wire [63:0] _GEN_2185 = write_counter[0] ? dcache_data_way0_1_rdata : dcache_data_way0_0_rdata; // @[data_cache.scala 356:{29,29}]
  wire  data_write_back_way = data_cache_under_write_back ? data_write_back_counter[7] : _GEN_384; // @[data_cache.scala 357:31]
  wire [63:0] writeback_data = data_write_back_way ? _GEN_2183 : _GEN_2185; // @[data_cache.scala 356:29]
  wire  _way0_burst_read_wen_T_2 = _wait_data_T_3 | _read_counter_T_9; // @[data_cache.scala 359:76]
  wire  _way0_burst_read_wen_T_4 = (_wait_data_T_3 | _read_counter_T_9) & io_port_rvalid; // @[data_cache.scala 359:124]
  wire  way0_burst_read_wen = (_wait_data_T_3 | _read_counter_T_9) & io_port_rvalid & _way0_dirty_T_7; // @[data_cache.scala 359:149]
  wire  way1_burst_read_wen = _way0_burst_read_wen_T_4 & _GEN_384; // @[data_cache.scala 360:149]
  wire  _dcache_data_way0_0_wdata_T_2 = _way0_dirty_T_9 | _way0_dirty_T; // @[data_cache.scala 363:81]
  wire [63:0] _dcache_data_way0_0_wdata_T_6 = _way0_burst_read_wen_T_2 ? io_port_rdata : 64'h0; // @[data_cache.scala 363:155]
  wire  _wen_way0_wire_0_T_1 = ~stage1_addr_line_mapping[3]; // @[data_cache.scala 373:59]
  wire  _way0_wen_0_T = 3'h0 == read_counter; // @[data_cache.scala 379:38]
  wire  way0_wen_0 = 3'h0 == read_counter & way0_burst_read_wen; // @[data_cache.scala 379:28]
  wire [7:0] _wen_way0_wire_0_T_13 = {way0_wen_0,way0_wen_0,way0_wen_0,way0_wen_0,way0_wen_0,way0_wen_0,way0_wen_0,
    way0_wen_0}; // @[Cat.scala 31:58]
  wire  way1_wen_0 = _way0_wen_0_T & way1_burst_read_wen; // @[data_cache.scala 380:28]
  wire [7:0] _wen_way1_wire_0_T_13 = {way1_wen_0,way1_wen_0,way1_wen_0,way1_wen_0,way1_wen_0,way1_wen_0,way1_wen_0,
    way1_wen_0}; // @[Cat.scala 31:58]
  wire  _way0_wen_1_T = 3'h1 == read_counter; // @[data_cache.scala 379:38]
  wire  way0_wen_1 = 3'h1 == read_counter & way0_burst_read_wen; // @[data_cache.scala 379:28]
  wire [7:0] _wen_way0_wire_1_T_13 = {way0_wen_1,way0_wen_1,way0_wen_1,way0_wen_1,way0_wen_1,way0_wen_1,way0_wen_1,
    way0_wen_1}; // @[Cat.scala 31:58]
  wire  way1_wen_1 = _way0_wen_1_T & way1_burst_read_wen; // @[data_cache.scala 380:28]
  wire [7:0] _wen_way1_wire_1_T_13 = {way1_wen_1,way1_wen_1,way1_wen_1,way1_wen_1,way1_wen_1,way1_wen_1,way1_wen_1,
    way1_wen_1}; // @[Cat.scala 31:58]
  wire [53:0] _T_27 = {1'h1,stage1_addr_line_mapping[63:11]}; // @[Cat.scala 31:58]
  wire  _io_port_araddr_T = work_state == 5'h1; // @[data_cache.scala 399:38]
  wire  _io_port_araddr_T_1 = work_state == 5'hc; // @[data_cache.scala 400:24]
  wire  _io_port_araddr_T_2 = work_state == 5'h8; // @[data_cache.scala 400:71]
  wire [63:0] _io_port_araddr_T_5 = {stage1_sram_phy_addr_reg[63:4],4'h0}; // @[Cat.scala 31:58]
  wire [63:0] _io_port_araddr_T_6 = work_state == 5'hc | work_state == 5'h8 ? _io_port_araddr_T_5 : 64'h0; // @[data_cache.scala 400:12]
  wire [1:0] _io_port_arsize_T_1 = stage1_sram_cache_reg ? 2'h3 : stage1_sram_size_reg; // @[data_cache.scala 402:27]
  wire  stage2_addr_same_as_stage1 = stage2_sram_addr_reg == stage1_addr_line_mapping; // @[data_cache.scala 411:56]
  wire  stage2_write_stage1_read = stage2_sram_write_reg & ~stage1_sram_wr_reg; // @[data_cache.scala 412:58]
  wire  _T_35 = work_state == 5'h3; // @[data_cache.scala 413:21]
  wire  _GEN_3338 = io_port_bvalid ? 1'h0 : write_access_complete_reg; // @[data_cache.scala 415:39 416:35 418:35]
  wire [52:0] _awaddr_miss_addr_T_2 = _way0_dirty_T_7 ? dcache_tag_io_tag : dcache_tag_1_io_tag; // @[data_cache.scala 421:36]
  wire [63:0] awaddr_miss_addr = {_awaddr_miss_addr_T_2,stage1_sram_phy_addr_reg[10:4],4'h0}; // @[Cat.scala 31:58]
  wire  _io_port_arvalid_T_7 = ~(stage2_addr_same_as_stage1 & stage2_write_stage1_read & write_access_complete_reg); // @[data_cache.scala 424:53]
  wire [52:0] _io_port_awaddr_T_1 = data_write_back_way ? dcache_tag_1_io_tag : dcache_tag_io_tag; // @[data_cache.scala 432:46]
  wire [63:0] _io_port_awaddr_T_3 = {_io_port_awaddr_T_1,data_write_back_counter[6:0],4'h0}; // @[Cat.scala 31:58]
  wire [63:0] _io_port_awaddr_T_5 = 5'h3 == work_state ? stage1_sram_phy_addr_reg : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _io_port_awaddr_T_7 = 5'h9 == work_state ? awaddr_miss_addr : _io_port_awaddr_T_5; // @[Mux.scala 81:58]
  wire [63:0] _io_port_awaddr_T_9 = 5'hf == work_state ? awaddr_miss_addr : _io_port_awaddr_T_7; // @[Mux.scala 81:58]
  wire  _io_port_awlen_T_2 = stage1_sram_cache_reg | _data_cache_under_write_back_T_3; // @[data_cache.scala 433:57]
  wire [1:0] _io_port_awsize_T_3 = _io_port_awlen_T_2 ? 2'h3 : stage1_sram_size_reg; // @[data_cache.scala 434:27]
  wire  _io_port_awvalid_T_4 = _T_35 | _write_counter_T_10 | _write_counter_T_1; // @[data_cache.scala 442:110]
  wire  _io_port_wdata_T = work_state == 5'h4; // @[data_cache.scala 446:38]
  wire  _io_port_wdata_T_2 = work_state == 5'h4 | _T_35; // @[data_cache.scala 446:67]
  wire  _io_port_wdata_T_7 = _write_counter_T_2 | _write_counter_T_10; // @[data_cache.scala 446:217]
  wire  _io_port_wdata_T_9 = _io_port_wdata_T_7 | _write_counter_T_9; // @[data_cache.scala 447:49]
  wire  _io_port_wdata_T_13 = _io_port_wdata_T_9 | _data_cache_under_write_back_T_3 | _data_cache_under_write_back_T_5; // @[data_cache.scala 448:51]
  wire [63:0] _io_port_wdata_T_14 = _io_port_wdata_T_13 ? writeback_data : 64'h0; // @[data_cache.scala 446:135]
  wire [7:0] _io_port_wstrb_T_14 = _io_port_wdata_T_13 ? 8'hff : 8'h0; // @[data_cache.scala 449:131]
  wire  _io_port_wlast_T_7 = _write_counter_T | _write_counter_T_9; // @[data_cache.scala 452:176]
  wire  _io_port_wlast_T_11 = _io_port_wlast_T_7 | _data_cache_under_write_back_T_3 | _data_cache_under_write_back_T_5; // @[data_cache.scala 453:53]
  wire  _io_port_wlast_T_13 = _io_port_wlast_T_11 & _access_work_state_T_23; // @[data_cache.scala 454:9]
  wire  _io_port_wvalid_T_8 = _io_port_wdata_T_2 | _write_counter_T | _write_counter_T_1 | _write_counter_T_10; // @[data_cache.scala 455:190]
  reg [63:0] sram_rdata_reg; // @[data_cache.scala 462:33]
  reg  stage2_stall_reg; // @[data_cache.scala 464:35]
  wire [63:0] _io_sram_rdata_T_2 = _data_cache_under_write_all_back_T_1 ? hit_word : 64'h0; // @[data_cache.scala 466:92]
  wire [63:0] _io_sram_rdata_T_3 = _data_cache_under_write_all_back_T ? wait_data : _io_sram_rdata_T_2; // @[data_cache.scala 466:46]
  dcache_tag dcache_tag ( // @[data_cache.scala 60:30]
    .clock(dcache_tag_clock),
    .reset(dcache_tag_reset),
    .io_wen(dcache_tag_io_wen),
    .io_wdata(dcache_tag_io_wdata),
    .io_raddr(dcache_tag_io_raddr),
    .io_waddr(dcache_tag_io_waddr),
    .io_hit(dcache_tag_io_hit),
    .io_valid(dcache_tag_io_valid),
    .io_tag(dcache_tag_io_tag),
    .io_w_valid(dcache_tag_io_w_valid)
  );
  dcache_tag dcache_tag_1 ( // @[data_cache.scala 61:30]
    .clock(dcache_tag_1_clock),
    .reset(dcache_tag_1_reset),
    .io_wen(dcache_tag_1_io_wen),
    .io_wdata(dcache_tag_1_io_wdata),
    .io_raddr(dcache_tag_1_io_raddr),
    .io_waddr(dcache_tag_1_io_waddr),
    .io_hit(dcache_tag_1_io_hit),
    .io_valid(dcache_tag_1_io_valid),
    .io_tag(dcache_tag_1_io_tag),
    .io_w_valid(dcache_tag_1_io_w_valid)
  );
  dcache_data dcache_data ( // @[data_cache.scala 93:62]
    .clock(dcache_data_clock),
    .io_wen(dcache_data_io_wen),
    .io_addr(dcache_data_io_addr),
    .io_wdata(dcache_data_io_wdata),
    .io_rdata(dcache_data_io_rdata)
  );
  dcache_data dcache_data_1 ( // @[data_cache.scala 93:62]
    .clock(dcache_data_1_clock),
    .io_wen(dcache_data_1_io_wen),
    .io_addr(dcache_data_1_io_addr),
    .io_wdata(dcache_data_1_io_wdata),
    .io_rdata(dcache_data_1_io_rdata)
  );
  dcache_data dcache_data_2 ( // @[data_cache.scala 94:62]
    .clock(dcache_data_2_clock),
    .io_wen(dcache_data_2_io_wen),
    .io_addr(dcache_data_2_io_addr),
    .io_wdata(dcache_data_2_io_wdata),
    .io_rdata(dcache_data_2_io_rdata)
  );
  dcache_data dcache_data_3 ( // @[data_cache.scala 94:62]
    .clock(dcache_data_3_clock),
    .io_wen(dcache_data_3_io_wen),
    .io_addr(dcache_data_3_io_addr),
    .io_wdata(dcache_data_3_io_wdata),
    .io_rdata(dcache_data_3_io_rdata)
  );
  assign io_port_araddr = work_state == 5'h1 ? stage1_sram_phy_addr_reg : _io_port_araddr_T_6; // @[data_cache.scala 399:26]
  assign io_port_arlen = {{3'd0}, stage1_sram_cache_reg}; // @[data_cache.scala 401:20]
  assign io_port_arsize = {{1'd0}, _io_port_arsize_T_1}; // @[data_cache.scala 402:20]
  assign io_port_arburst = {{1'd0}, stage1_sram_cache_reg}; // @[data_cache.scala 406:21]
  assign io_port_arvalid = (_io_port_araddr_T | _io_port_araddr_T_1 | _io_port_araddr_T_2) & _io_port_arvalid_T_7; // @[data_cache.scala 423:27]
  assign io_port_awaddr = 5'h12 == work_state ? _io_port_awaddr_T_3 : _io_port_awaddr_T_9; // @[Mux.scala 81:58]
  assign io_port_awlen = {{3'd0}, _io_port_awlen_T_2}; // @[data_cache.scala 433:21]
  assign io_port_awsize = {{1'd0}, _io_port_awsize_T_3}; // @[data_cache.scala 434:21]
  assign io_port_awburst = {{1'd0}, _io_port_awlen_T_2}; // @[data_cache.scala 438:21]
  assign io_port_awvalid = _io_port_awvalid_T_4 | _data_cache_under_write_back_T_3; // @[data_cache.scala 443:10]
  assign io_port_wdata = work_state == 5'h4 | _T_35 ? stage1_sram_wdata_reg : _io_port_wdata_T_14; // @[data_cache.scala 446:26]
  assign io_port_wstrb = _io_port_wdata_T_2 ? stage1_wstrb_reg : _io_port_wstrb_T_14; // @[data_cache.scala 449:26]
  assign io_port_wlast = _io_port_wdata_T | _T_35 & io_port_wready | _io_port_wlast_T_13; // @[data_cache.scala 452:132]
  assign io_port_wvalid = _io_port_wvalid_T_8 | _write_counter_T_9 | _data_cache_under_write_back_T_3 |
    _data_cache_under_write_back_T_5; // @[data_cache.scala 456:136]
  assign io_stage2_stall = access_work_state_for_stall[4:3] == 2'h3; // @[data_cache.scala 288:54]
  assign io_v_addr_for_tlb = stage1_addr_line_mapping; // @[data_cache.scala 222:23]
  assign io_tlb_req = _io_tlb_req_T_4 & stage1_sram_req_reg; // @[data_cache.scala 221:54]
  assign io_sram_rdata = stage2_stall_reg ? _io_sram_rdata_T_3 : sram_rdata_reg; // @[data_cache.scala 466:25]
  assign dcache_tag_clock = clock;
  assign dcache_tag_reset = reset;
  assign dcache_tag_io_wen = _way0_burst_read_wen_T_2 & _way0_dirty_T_7; // @[data_cache.scala 389:122]
  assign dcache_tag_io_wdata = _way0_burst_read_wen_T_2 ? _T_27 : 54'h0; // @[data_cache.scala 391:30]
  assign dcache_tag_io_raddr = io_sram_addr; // @[data_cache.scala 216:24]
  assign dcache_tag_io_waddr = data_cache_under_write_back ? {{53'd0}, _T_3} : stage1_addr_line_mapping; // @[data_cache.scala 213:30]
  assign dcache_tag_1_clock = clock;
  assign dcache_tag_1_reset = reset;
  assign dcache_tag_1_io_wen = _way0_burst_read_wen_T_2 & _GEN_384; // @[data_cache.scala 390:122]
  assign dcache_tag_1_io_wdata = _way0_burst_read_wen_T_2 ? _T_27 : 54'h0; // @[data_cache.scala 392:30]
  assign dcache_tag_1_io_raddr = io_sram_addr; // @[data_cache.scala 217:24]
  assign dcache_tag_1_io_waddr = data_cache_under_write_back ? {{53'd0}, _T_3} : stage1_addr_line_mapping; // @[data_cache.scala 214:30]
  assign dcache_data_clock = clock;
  assign dcache_data_io_wen = ~stage1_addr_line_mapping[3] & (_way0_dirty_T_4 | _way0_dirty_T_12) ? stage1_wstrb_reg :
    _wen_way0_wire_0_T_13; // @[data_cache.scala 373:33]
  assign dcache_data_io_addr = data_cache_under_write_back ? {{53'd0}, _T_3} : stage1_addr_line_mapping; // @[data_cache.scala 362:40]
  assign dcache_data_io_wdata = _way0_dirty_T_9 | _way0_dirty_T ? stage1_sram_wdata_reg : _dcache_data_way0_0_wdata_T_6; // @[data_cache.scala 363:41]
  assign dcache_data_1_clock = clock;
  assign dcache_data_1_io_wen = stage1_addr_line_mapping[3] & (_way0_dirty_T_4 | _way0_dirty_T_12) ? stage1_wstrb_reg :
    _wen_way0_wire_1_T_13; // @[data_cache.scala 373:33]
  assign dcache_data_1_io_addr = data_cache_under_write_back ? {{53'd0}, _T_3} : stage1_addr_line_mapping; // @[data_cache.scala 362:40]
  assign dcache_data_1_io_wdata = _way0_dirty_T_9 | _way0_dirty_T ? stage1_sram_wdata_reg :
    _dcache_data_way0_0_wdata_T_6; // @[data_cache.scala 363:41]
  assign dcache_data_2_clock = clock;
  assign dcache_data_2_io_wen = _wen_way0_wire_0_T_1 & (_way1_dirty_T_4 | _way1_dirty_T_12) ? stage1_wstrb_reg :
    _wen_way1_wire_0_T_13; // @[data_cache.scala 375:33]
  assign dcache_data_2_io_addr = data_cache_under_write_back ? {{53'd0}, _T_3} : stage1_addr_line_mapping; // @[data_cache.scala 366:40]
  assign dcache_data_2_io_wdata = _dcache_data_way0_0_wdata_T_2 ? stage1_sram_wdata_reg : _dcache_data_way0_0_wdata_T_6; // @[data_cache.scala 367:41]
  assign dcache_data_3_clock = clock;
  assign dcache_data_3_io_wen = stage1_addr_line_mapping[3] & (_way1_dirty_T_4 | _way1_dirty_T_12) ? stage1_wstrb_reg :
    _wen_way1_wire_1_T_13; // @[data_cache.scala 375:33]
  assign dcache_data_3_io_addr = data_cache_under_write_back ? {{53'd0}, _T_3} : stage1_addr_line_mapping; // @[data_cache.scala 366:40]
  assign dcache_data_3_io_wdata = _dcache_data_way0_0_wdata_T_2 ? stage1_sram_wdata_reg : _dcache_data_way0_0_wdata_T_6; // @[data_cache.scala 367:41]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Mux.scala 81:58]
      work_state <= 5'h18; // @[data_cache.scala 274:41]
    end else if (5'h15 == work_state) begin // @[Mux.scala 81:58]
      if (data_all_write_back) begin // @[data_cache.scala 273:41]
        work_state <= 5'h18;
      end else begin
        work_state <= 5'h11;
      end
    end else if (5'h14 == work_state) begin // @[Mux.scala 81:58]
      if (io_port_bvalid) begin // @[data_cache.scala 272:41]
        work_state <= 5'h15;
      end
    end else if (5'h13 == work_state) begin // @[Mux.scala 81:58]
      if (_access_work_state_T_24) begin
        work_state <= 5'h14;
      end
    end else if (5'h12 == work_state) begin
      work_state <= _access_work_state_T_45;
    end else begin
      work_state <= _access_work_state_T_92;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 295:25]
      write_counter <= 3'h0;
    end else if (work_state == 5'ha | work_state == 5'h9) begin // @[data_cache.scala 296:12]
      write_counter <= _write_counter_T_8;
    end else if (work_state == 5'h6 | work_state == 5'hf) begin // @[data_cache.scala 297:12]
      write_counter <= _write_counter_T_8;
    end else if (_data_cache_under_write_back_T_5 | _data_cache_under_write_back_T_3) begin
      write_counter <= _write_counter_T_8;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 298:24]
      read_counter <= 3'h0;
    end else if (_wait_data_T_3) begin // @[data_cache.scala 299:12]
      read_counter <= _read_counter_T_8;
    end else if (work_state == 5'h0) begin
      read_counter <= _read_counter_T_8;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 292:21]
      wait_data <= 64'h0;
    end else if (work_state == 5'h2 & io_port_rvalid) begin // @[data_cache.scala 293:12]
      wait_data <= io_port_rdata;
    end else if (work_state == 5'hd & io_port_rvalid & read_counter == _GEN_3468) begin
      wait_data <= io_port_rdata;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_0 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h0 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_0 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_0 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_0 <= lru_127;
      end else begin
        lru_0 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_1 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h1 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_1 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_1 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_1 <= lru_127;
      end else begin
        lru_1 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_2 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h2 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_2 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_2 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_2 <= lru_127;
      end else begin
        lru_2 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_3 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h3 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_3 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_3 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_3 <= lru_127;
      end else begin
        lru_3 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_4 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h4 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_4 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_4 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_4 <= lru_127;
      end else begin
        lru_4 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_5 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h5 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_5 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_5 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_5 <= lru_127;
      end else begin
        lru_5 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_6 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h6 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_6 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_6 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_6 <= lru_127;
      end else begin
        lru_6 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_7 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h7 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_7 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_7 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_7 <= lru_127;
      end else begin
        lru_7 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_8 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h8 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_8 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_8 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_8 <= lru_127;
      end else begin
        lru_8 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_9 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h9 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_9 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_9 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_9 <= lru_127;
      end else begin
        lru_9 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_10 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'ha == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_10 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_10 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_10 <= lru_127;
      end else begin
        lru_10 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_11 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'hb == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_11 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_11 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_11 <= lru_127;
      end else begin
        lru_11 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_12 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'hc == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_12 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_12 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_12 <= lru_127;
      end else begin
        lru_12 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_13 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'hd == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_13 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_13 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_13 <= lru_127;
      end else begin
        lru_13 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_14 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'he == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_14 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_14 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_14 <= lru_127;
      end else begin
        lru_14 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_15 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'hf == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_15 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_15 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_15 <= lru_127;
      end else begin
        lru_15 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_16 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h10 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_16 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_16 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_16 <= lru_127;
      end else begin
        lru_16 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_17 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h11 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_17 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_17 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_17 <= lru_127;
      end else begin
        lru_17 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_18 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h12 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_18 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_18 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_18 <= lru_127;
      end else begin
        lru_18 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_19 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h13 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_19 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_19 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_19 <= lru_127;
      end else begin
        lru_19 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_20 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h14 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_20 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_20 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_20 <= lru_127;
      end else begin
        lru_20 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_21 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h15 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_21 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_21 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_21 <= lru_127;
      end else begin
        lru_21 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_22 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h16 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_22 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_22 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_22 <= lru_127;
      end else begin
        lru_22 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_23 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h17 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_23 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_23 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_23 <= lru_127;
      end else begin
        lru_23 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_24 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h18 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_24 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_24 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_24 <= lru_127;
      end else begin
        lru_24 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_25 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h19 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_25 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_25 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_25 <= lru_127;
      end else begin
        lru_25 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_26 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h1a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_26 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_26 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_26 <= lru_127;
      end else begin
        lru_26 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_27 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h1b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_27 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_27 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_27 <= lru_127;
      end else begin
        lru_27 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_28 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h1c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_28 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_28 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_28 <= lru_127;
      end else begin
        lru_28 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_29 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h1d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_29 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_29 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_29 <= lru_127;
      end else begin
        lru_29 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_30 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h1e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_30 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_30 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_30 <= lru_127;
      end else begin
        lru_30 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_31 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h1f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_31 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_31 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_31 <= lru_127;
      end else begin
        lru_31 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_32 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h20 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_32 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_32 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_32 <= lru_127;
      end else begin
        lru_32 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_33 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h21 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_33 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_33 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_33 <= lru_127;
      end else begin
        lru_33 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_34 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h22 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_34 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_34 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_34 <= lru_127;
      end else begin
        lru_34 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_35 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h23 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_35 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_35 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_35 <= lru_127;
      end else begin
        lru_35 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_36 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h24 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_36 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_36 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_36 <= lru_127;
      end else begin
        lru_36 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_37 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h25 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_37 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_37 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_37 <= lru_127;
      end else begin
        lru_37 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_38 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h26 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_38 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_38 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_38 <= lru_127;
      end else begin
        lru_38 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_39 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h27 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_39 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_39 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_39 <= lru_127;
      end else begin
        lru_39 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_40 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h28 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_40 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_40 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_40 <= lru_127;
      end else begin
        lru_40 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_41 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h29 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_41 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_41 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_41 <= lru_127;
      end else begin
        lru_41 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_42 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h2a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_42 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_42 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_42 <= lru_127;
      end else begin
        lru_42 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_43 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h2b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_43 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_43 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_43 <= lru_127;
      end else begin
        lru_43 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_44 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h2c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_44 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_44 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_44 <= lru_127;
      end else begin
        lru_44 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_45 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h2d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_45 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_45 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_45 <= lru_127;
      end else begin
        lru_45 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_46 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h2e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_46 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_46 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_46 <= lru_127;
      end else begin
        lru_46 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_47 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h2f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_47 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_47 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_47 <= lru_127;
      end else begin
        lru_47 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_48 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h30 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_48 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_48 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_48 <= lru_127;
      end else begin
        lru_48 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_49 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h31 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_49 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_49 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_49 <= lru_127;
      end else begin
        lru_49 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_50 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h32 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_50 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_50 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_50 <= lru_127;
      end else begin
        lru_50 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_51 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h33 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_51 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_51 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_51 <= lru_127;
      end else begin
        lru_51 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_52 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h34 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_52 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_52 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_52 <= lru_127;
      end else begin
        lru_52 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_53 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h35 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_53 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_53 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_53 <= lru_127;
      end else begin
        lru_53 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_54 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h36 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_54 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_54 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_54 <= lru_127;
      end else begin
        lru_54 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_55 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h37 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_55 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_55 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_55 <= lru_127;
      end else begin
        lru_55 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_56 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h38 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_56 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_56 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_56 <= lru_127;
      end else begin
        lru_56 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_57 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h39 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_57 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_57 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_57 <= lru_127;
      end else begin
        lru_57 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_58 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h3a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_58 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_58 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_58 <= lru_127;
      end else begin
        lru_58 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_59 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h3b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_59 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_59 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_59 <= lru_127;
      end else begin
        lru_59 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_60 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h3c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_60 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_60 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_60 <= lru_127;
      end else begin
        lru_60 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_61 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h3d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_61 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_61 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_61 <= lru_127;
      end else begin
        lru_61 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_62 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h3e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_62 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_62 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_62 <= lru_127;
      end else begin
        lru_62 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_63 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h3f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_63 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_63 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_63 <= lru_127;
      end else begin
        lru_63 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_64 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h40 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_64 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_64 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_64 <= lru_127;
      end else begin
        lru_64 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_65 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h41 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_65 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_65 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_65 <= lru_127;
      end else begin
        lru_65 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_66 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h42 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_66 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_66 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_66 <= lru_127;
      end else begin
        lru_66 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_67 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h43 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_67 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_67 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_67 <= lru_127;
      end else begin
        lru_67 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_68 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h44 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_68 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_68 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_68 <= lru_127;
      end else begin
        lru_68 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_69 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h45 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_69 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_69 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_69 <= lru_127;
      end else begin
        lru_69 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_70 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h46 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_70 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_70 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_70 <= lru_127;
      end else begin
        lru_70 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_71 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h47 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_71 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_71 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_71 <= lru_127;
      end else begin
        lru_71 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_72 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h48 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_72 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_72 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_72 <= lru_127;
      end else begin
        lru_72 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_73 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h49 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_73 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_73 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_73 <= lru_127;
      end else begin
        lru_73 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_74 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h4a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_74 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_74 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_74 <= lru_127;
      end else begin
        lru_74 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_75 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h4b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_75 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_75 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_75 <= lru_127;
      end else begin
        lru_75 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_76 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h4c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_76 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_76 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_76 <= lru_127;
      end else begin
        lru_76 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_77 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h4d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_77 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_77 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_77 <= lru_127;
      end else begin
        lru_77 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_78 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h4e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_78 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_78 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_78 <= lru_127;
      end else begin
        lru_78 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_79 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h4f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_79 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_79 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_79 <= lru_127;
      end else begin
        lru_79 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_80 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h50 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_80 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_80 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_80 <= lru_127;
      end else begin
        lru_80 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_81 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h51 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_81 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_81 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_81 <= lru_127;
      end else begin
        lru_81 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_82 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h52 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_82 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_82 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_82 <= lru_127;
      end else begin
        lru_82 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_83 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h53 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_83 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_83 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_83 <= lru_127;
      end else begin
        lru_83 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_84 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h54 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_84 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_84 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_84 <= lru_127;
      end else begin
        lru_84 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_85 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h55 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_85 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_85 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_85 <= lru_127;
      end else begin
        lru_85 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_86 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h56 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_86 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_86 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_86 <= lru_127;
      end else begin
        lru_86 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_87 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h57 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_87 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_87 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_87 <= lru_127;
      end else begin
        lru_87 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_88 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h58 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_88 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_88 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_88 <= lru_127;
      end else begin
        lru_88 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_89 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h59 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_89 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_89 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_89 <= lru_127;
      end else begin
        lru_89 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_90 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h5a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_90 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_90 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_90 <= lru_127;
      end else begin
        lru_90 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_91 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h5b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_91 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_91 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_91 <= lru_127;
      end else begin
        lru_91 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_92 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h5c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_92 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_92 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_92 <= lru_127;
      end else begin
        lru_92 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_93 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h5d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_93 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_93 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_93 <= lru_127;
      end else begin
        lru_93 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_94 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h5e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_94 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_94 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_94 <= lru_127;
      end else begin
        lru_94 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_95 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h5f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_95 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_95 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_95 <= lru_127;
      end else begin
        lru_95 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_96 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h60 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_96 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_96 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_96 <= lru_127;
      end else begin
        lru_96 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_97 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h61 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_97 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_97 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_97 <= lru_127;
      end else begin
        lru_97 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_98 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h62 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_98 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_98 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_98 <= lru_127;
      end else begin
        lru_98 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_99 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h63 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_99 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_99 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_99 <= lru_127;
      end else begin
        lru_99 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_100 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h64 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_100 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_100 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_100 <= lru_127;
      end else begin
        lru_100 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_101 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h65 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_101 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_101 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_101 <= lru_127;
      end else begin
        lru_101 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_102 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h66 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_102 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_102 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_102 <= lru_127;
      end else begin
        lru_102 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_103 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h67 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_103 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_103 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_103 <= lru_127;
      end else begin
        lru_103 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_104 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h68 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_104 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_104 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_104 <= lru_127;
      end else begin
        lru_104 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_105 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h69 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_105 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_105 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_105 <= lru_127;
      end else begin
        lru_105 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_106 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h6a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_106 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_106 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_106 <= lru_127;
      end else begin
        lru_106 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_107 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h6b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_107 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_107 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_107 <= lru_127;
      end else begin
        lru_107 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_108 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h6c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_108 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_108 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_108 <= lru_127;
      end else begin
        lru_108 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_109 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h6d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_109 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_109 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_109 <= lru_127;
      end else begin
        lru_109 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_110 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h6e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_110 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_110 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_110 <= lru_127;
      end else begin
        lru_110 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_111 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h6f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_111 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_111 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_111 <= lru_127;
      end else begin
        lru_111 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_112 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h70 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_112 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_112 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_112 <= lru_127;
      end else begin
        lru_112 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_113 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h71 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_113 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_113 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_113 <= lru_127;
      end else begin
        lru_113 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_114 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h72 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_114 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_114 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_114 <= lru_127;
      end else begin
        lru_114 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_115 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h73 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_115 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_115 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_115 <= lru_127;
      end else begin
        lru_115 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_116 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h74 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_116 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_116 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_116 <= lru_127;
      end else begin
        lru_116 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_117 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h75 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_117 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_117 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_117 <= lru_127;
      end else begin
        lru_117 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_118 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h76 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_118 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_118 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_118 <= lru_127;
      end else begin
        lru_118 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_119 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h77 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_119 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_119 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_119 <= lru_127;
      end else begin
        lru_119 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_120 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h78 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_120 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_120 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_120 <= lru_127;
      end else begin
        lru_120 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_121 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h79 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_121 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_121 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_121 <= lru_127;
      end else begin
        lru_121 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_122 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h7a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_122 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_122 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_122 <= lru_127;
      end else begin
        lru_122 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_123 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h7b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_123 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_123 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_123 <= lru_127;
      end else begin
        lru_123 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_124 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h7c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_124 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_124 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_124 <= lru_127;
      end else begin
        lru_124 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_125 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h7d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_125 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_125 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_125 <= lru_127;
      end else begin
        lru_125 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_126 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h7e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_126 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_126 <= _way0_dirty_T_7;
      end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin
        lru_126 <= lru_127;
      end else begin
        lru_126 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 228:37]
      lru_127 <= 1'h0; // @[data_cache.scala 228:43 231:12 200:{86,86}]
    end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 63:22]
      if (_way0_dirty_T) begin
        lru_127 <= _lru_T_5;
      end else if (_way0_dirty_T_5 | _way0_dirty_T_9) begin
        lru_127 <= _way0_dirty_T_7;
      end else if (!(7'h7f == stage1_addr_line_mapping[10:4])) begin
        lru_127 <= _GEN_383;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_0 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h0 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_0 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_1 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h1 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_1 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_2 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h2 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_2 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_3 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h3 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_3 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_4 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h4 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_4 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_5 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h5 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_5 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_6 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h6 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_6 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_7 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h7 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_7 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_8 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h8 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_8 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_9 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h9 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_9 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_10 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'ha == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_10 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_11 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'hb == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_11 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_12 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'hc == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_12 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_13 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'hd == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_13 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_14 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'he == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_14 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_15 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'hf == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_15 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_16 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h10 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_16 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_17 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h11 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_17 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_18 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h12 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_18 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_19 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h13 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_19 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_20 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h14 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_20 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_21 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h15 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_21 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_22 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h16 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_22 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_23 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h17 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_23 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_24 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h18 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_24 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_25 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h19 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_25 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_26 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h1a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_26 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_27 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h1b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_27 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_28 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h1c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_28 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_29 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h1d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_29 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_30 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h1e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_30 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_31 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h1f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_31 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_32 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h20 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_32 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_33 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h21 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_33 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_34 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h22 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_34 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_35 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h23 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_35 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_36 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h24 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_36 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_37 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h25 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_37 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_38 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h26 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_38 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_39 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h27 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_39 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_40 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h28 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_40 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_41 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h29 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_41 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_42 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h2a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_42 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_43 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h2b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_43 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_44 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h2c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_44 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_45 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h2d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_45 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_46 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h2e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_46 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_47 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h2f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_47 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_48 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h30 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_48 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_49 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h31 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_49 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_50 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h32 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_50 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_51 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h33 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_51 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_52 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h34 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_52 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_53 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h35 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_53 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_54 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h36 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_54 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_55 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h37 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_55 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_56 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h38 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_56 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_57 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h39 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_57 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_58 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h3a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_58 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_59 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h3b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_59 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_60 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h3c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_60 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_61 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h3d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_61 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_62 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h3e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_62 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_63 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h3f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_63 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_64 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h40 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_64 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_65 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h41 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_65 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_66 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h42 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_66 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_67 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h43 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_67 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_68 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h44 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_68 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_69 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h45 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_69 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_70 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h46 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_70 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_71 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h47 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_71 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_72 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h48 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_72 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_73 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h49 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_73 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_74 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h4a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_74 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_75 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h4b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_75 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_76 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h4c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_76 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_77 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h4d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_77 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_78 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h4e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_78 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_79 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h4f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_79 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_80 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h50 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_80 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_81 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h51 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_81 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_82 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h52 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_82 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_83 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h53 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_83 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_84 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h54 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_84 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_85 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h55 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_85 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_86 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h56 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_86 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_87 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h57 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_87 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_88 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h58 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_88 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_89 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h59 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_89 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_90 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h5a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_90 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_91 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h5b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_91 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_92 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h5c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_92 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_93 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h5d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_93 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_94 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h5e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_94 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_95 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h5f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_95 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_96 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h60 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_96 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_97 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h61 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_97 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_98 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h62 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_98 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_99 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h63 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_99 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_100 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h64 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_100 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_101 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h65 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_101 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_102 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h66 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_102 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_103 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h67 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_103 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_104 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h68 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_104 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_105 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h69 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_105 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_106 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h6a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_106 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_107 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h6b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_107 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_108 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h6c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_108 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_109 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h6d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_109 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_110 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h6e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_110 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_111 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h6f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_111 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_112 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h70 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_112 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_113 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h71 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_113 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_114 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h72 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_114 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_115 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h73 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_115 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_116 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h74 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_116 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_117 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h75 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_117 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_118 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h76 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_118 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_119 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h77 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_119 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_120 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h78 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_120 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_121 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h79 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_121 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_122 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h7a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_122 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_123 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h7b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_123 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_124 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h7c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_124 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_125 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h7d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_125 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_126 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h7e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_126 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 199:44]
      way0_dirty_127 <= 1'h0; // @[data_cache.scala 199:44]
    end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 64:29]
      way0_dirty_127 <= state_lookup_for_less_delay == 5'h19 & stage1_sram_wr_reg & stage1_sram_hit0_reg &
        stage1_sram_valid0_reg | _way0_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_0 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h0 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_0 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_1 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h1 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_1 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_2 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h2 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_2 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_3 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h3 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_3 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_4 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h4 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_4 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_5 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h5 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_5 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_6 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h6 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_6 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_7 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h7 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_7 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_8 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h8 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_8 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_9 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h9 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_9 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_10 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'ha == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_10 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_11 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'hb == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_11 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_12 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'hc == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_12 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_13 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'hd == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_13 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_14 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'he == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_14 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_15 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'hf == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_15 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_16 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h10 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_16 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_17 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h11 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_17 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_18 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h12 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_18 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_19 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h13 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_19 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_20 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h14 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_20 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_21 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h15 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_21 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_22 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h16 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_22 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_23 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h17 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_23 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_24 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h18 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_24 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_25 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h19 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_25 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_26 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h1a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_26 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_27 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h1b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_27 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_28 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h1c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_28 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_29 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h1d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_29 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_30 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h1e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_30 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_31 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h1f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_31 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_32 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h20 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_32 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_33 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h21 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_33 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_34 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h22 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_34 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_35 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h23 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_35 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_36 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h24 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_36 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_37 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h25 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_37 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_38 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h26 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_38 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_39 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h27 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_39 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_40 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h28 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_40 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_41 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h29 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_41 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_42 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h2a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_42 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_43 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h2b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_43 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_44 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h2c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_44 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_45 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h2d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_45 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_46 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h2e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_46 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_47 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h2f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_47 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_48 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h30 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_48 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_49 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h31 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_49 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_50 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h32 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_50 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_51 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h33 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_51 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_52 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h34 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_52 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_53 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h35 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_53 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_54 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h36 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_54 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_55 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h37 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_55 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_56 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h38 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_56 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_57 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h39 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_57 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_58 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h3a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_58 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_59 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h3b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_59 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_60 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h3c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_60 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_61 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h3d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_61 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_62 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h3e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_62 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_63 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h3f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_63 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_64 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h40 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_64 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_65 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h41 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_65 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_66 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h42 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_66 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_67 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h43 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_67 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_68 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h44 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_68 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_69 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h45 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_69 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_70 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h46 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_70 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_71 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h47 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_71 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_72 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h48 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_72 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_73 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h49 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_73 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_74 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h4a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_74 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_75 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h4b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_75 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_76 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h4c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_76 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_77 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h4d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_77 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_78 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h4e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_78 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_79 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h4f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_79 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_80 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h50 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_80 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_81 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h51 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_81 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_82 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h52 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_82 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_83 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h53 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_83 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_84 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h54 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_84 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_85 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h55 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_85 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_86 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h56 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_86 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_87 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h57 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_87 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_88 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h58 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_88 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_89 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h59 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_89 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_90 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h5a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_90 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_91 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h5b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_91 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_92 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h5c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_92 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_93 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h5d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_93 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_94 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h5e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_94 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_95 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h5f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_95 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_96 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h60 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_96 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_97 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h61 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_97 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_98 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h62 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_98 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_99 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h63 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_99 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_100 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h64 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_100 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_101 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h65 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_101 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_102 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h66 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_102 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_103 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h67 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_103 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_104 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h68 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_104 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_105 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h69 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_105 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_106 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h6a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_106 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_107 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h6b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_107 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_108 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h6c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_108 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_109 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h6d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_109 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_110 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h6e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_110 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_111 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h6f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_111 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_112 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h70 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_112 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_113 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h71 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_113 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_114 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h72 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_114 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_115 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h73 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_115 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_116 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h74 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_116 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_117 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h75 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_117 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_118 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h76 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_118 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_119 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h77 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_119 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_120 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h78 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_120 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_121 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h79 == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_121 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_122 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h7a == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_122 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_123 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h7b == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_123 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_124 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h7c == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_124 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_125 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h7d == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_125 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_126 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h7e == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_126 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 203:44]
      way1_dirty_127 <= 1'h0; // @[data_cache.scala 203:44]
    end else if (7'h7f == stage1_addr_line_mapping[10:4]) begin // @[data_cache.scala 65:29]
      way1_dirty_127 <= _way0_dirty_T_2 & stage1_sram_hit1_reg & stage1_sram_valid1_reg | _way1_dirty_T_15;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 185:32]
      stage1_addr_line_mapping <= 64'h0;
    end else if (io_sram_req) begin
      stage1_addr_line_mapping <= io_sram_addr;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 186:33]
      stage1_sram_cache_reg <= 1'h0;
    end else if (io_sram_req) begin
      stage1_sram_cache_reg <= io_sram_cache;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 187:33]
      stage1_sram_wdata_reg <= 64'h0;
    end else if (io_sram_req) begin
      stage1_sram_wdata_reg <= io_sram_wdata;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 72:39]
      stage1_sram_size_reg <= 2'h0; // @[data_cache.scala 72:39]
    end else begin
      stage1_sram_size_reg <= _stage1_sram_size_reg_T_1[1:0]; // @[data_cache.scala 188:27]
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 189:33]
      stage1_sram_wr_reg <= 1'h0;
    end else if (io_sram_req) begin
      stage1_sram_wr_reg <= io_sram_wr;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 190:33]
      stage1_sram_req_reg <= 1'h0;
    end else begin
      stage1_sram_req_reg <= io_sram_req | _stage1_sram_req_reg_T_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 193:32]
      stage1_sram_hit0_reg <= 1'h0;
    end else if (io_sram_req) begin
      stage1_sram_hit0_reg <= dcache_tag_io_hit;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 194:32]
      stage1_sram_hit1_reg <= 1'h0;
    end else if (io_sram_req) begin
      stage1_sram_hit1_reg <= dcache_tag_1_io_hit;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 195:34]
      stage1_sram_valid0_reg <= 1'h0;
    end else if (io_sram_req) begin
      stage1_sram_valid0_reg <= dcache_tag_io_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 196:34]
      stage1_sram_valid1_reg <= 1'h0;
    end else if (io_sram_req) begin
      stage1_sram_valid1_reg <= dcache_tag_1_io_valid;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 191:33]
      stage1_wstrb_reg <= 8'h0;
    end else if (io_sram_req) begin
      stage1_wstrb_reg <= io_data_wstrb;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 224:37]
      stage1_sram_phy_addr_reg <= 64'h0; // @[data_cache.scala 224:73]
    end else if (stage1_stall_reg) begin
      if (io_tlb_req) begin
        stage1_sram_phy_addr_reg <= io_p_addr_for_tlb;
      end else begin
        stage1_sram_phy_addr_reg <= stage1_addr_line_mapping;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Mux.scala 101:16]
      data_write_back_counter <= 8'h0;
    end else if (_data_write_back_counter_T_2) begin // @[Mux.scala 101:16]
      data_write_back_counter <= _data_write_back_counter_T_4;
    end else if (_data_cache_under_write_back_T_1) begin
      data_write_back_counter <= _data_write_back_counter_T_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 318:54]
      stage2_sram_write_reg <= 1'h0;
    end else if (stage2_stall) begin
      stage2_sram_write_reg <= stage1_sram_wr_reg;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 179:37]
      stage1_stall_reg <= 1'h0;
    end else begin
      stage1_stall_reg <= io_sram_req;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 413:52]
      write_access_complete_reg <= 1'h0; // @[data_cache.scala 414:35]
    end else begin
      write_access_complete_reg <= work_state == 5'h3 | _GEN_3338;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Reg.scala 29:18]
      stage2_sram_addr_reg <= 64'h0; // @[Reg.scala 29:22]
    end else if (stage2_stall) begin // @[Reg.scala 28:20]
      stage2_sram_addr_reg <= stage1_addr_line_mapping;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 322:48]
      stage2_hit0_reg <= 1'h0;
    end else if (stage2_stall) begin
      stage2_hit0_reg <= _hit_T;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 463:27]
      sram_rdata_reg <= 64'h0;
    end else if (_data_cache_under_write_all_back_T) begin // @[data_cache.scala 463:73]
      sram_rdata_reg <= wait_data; // @[data_cache.scala 346:{23,23,23,23,23}]
    end else if (_data_cache_under_write_all_back_T_1) begin
      if (stage2_hit0_reg) begin
        if (stage2_sram_addr_reg[3]) begin
          sram_rdata_reg <= dcache_data_way0_1_rdata;
        end else begin
          sram_rdata_reg <= dcache_data_way0_0_rdata;
        end
      end else if (stage2_sram_addr_reg[3]) begin
        sram_rdata_reg <= dcache_data_way1_1_rdata;
      end else begin
        sram_rdata_reg <= dcache_data_way1_0_rdata;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[data_cache.scala 288:54]
      stage2_stall_reg <= 1'h0;
    end else begin
      stage2_stall_reg <= access_work_state_for_stall[4:3] == 2'h3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  work_state = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  write_counter = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  read_counter = _RAND_2[2:0];
  _RAND_3 = {2{`RANDOM}};
  wait_data = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  lru_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lru_1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  lru_2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  lru_3 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  lru_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  lru_5 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  lru_6 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  lru_7 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  lru_8 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  lru_9 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  lru_10 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  lru_11 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  lru_12 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  lru_13 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  lru_14 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  lru_15 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  lru_16 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  lru_17 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  lru_18 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  lru_19 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  lru_20 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  lru_21 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  lru_22 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  lru_23 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  lru_24 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  lru_25 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  lru_26 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  lru_27 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  lru_28 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  lru_29 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  lru_30 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  lru_31 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  lru_32 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  lru_33 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  lru_34 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  lru_35 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  lru_36 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  lru_37 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  lru_38 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  lru_39 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  lru_40 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  lru_41 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  lru_42 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  lru_43 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  lru_44 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  lru_45 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  lru_46 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  lru_47 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  lru_48 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  lru_49 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  lru_50 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  lru_51 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  lru_52 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  lru_53 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  lru_54 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  lru_55 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  lru_56 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  lru_57 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  lru_58 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  lru_59 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  lru_60 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  lru_61 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  lru_62 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  lru_63 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  lru_64 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  lru_65 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  lru_66 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  lru_67 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  lru_68 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  lru_69 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  lru_70 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  lru_71 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  lru_72 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  lru_73 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  lru_74 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  lru_75 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  lru_76 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  lru_77 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  lru_78 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  lru_79 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  lru_80 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  lru_81 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  lru_82 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  lru_83 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  lru_84 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  lru_85 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  lru_86 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  lru_87 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  lru_88 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  lru_89 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  lru_90 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  lru_91 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  lru_92 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  lru_93 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  lru_94 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  lru_95 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  lru_96 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  lru_97 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  lru_98 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  lru_99 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  lru_100 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  lru_101 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  lru_102 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  lru_103 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  lru_104 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  lru_105 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  lru_106 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  lru_107 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  lru_108 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  lru_109 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  lru_110 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  lru_111 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  lru_112 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  lru_113 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  lru_114 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  lru_115 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  lru_116 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  lru_117 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  lru_118 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  lru_119 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  lru_120 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  lru_121 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  lru_122 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  lru_123 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  lru_124 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  lru_125 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  lru_126 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  lru_127 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  way0_dirty_0 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  way0_dirty_1 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  way0_dirty_2 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  way0_dirty_3 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  way0_dirty_4 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  way0_dirty_5 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  way0_dirty_6 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  way0_dirty_7 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  way0_dirty_8 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  way0_dirty_9 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  way0_dirty_10 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  way0_dirty_11 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  way0_dirty_12 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  way0_dirty_13 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  way0_dirty_14 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  way0_dirty_15 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  way0_dirty_16 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  way0_dirty_17 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  way0_dirty_18 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  way0_dirty_19 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  way0_dirty_20 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  way0_dirty_21 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  way0_dirty_22 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  way0_dirty_23 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  way0_dirty_24 = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  way0_dirty_25 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  way0_dirty_26 = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  way0_dirty_27 = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  way0_dirty_28 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  way0_dirty_29 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  way0_dirty_30 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  way0_dirty_31 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  way0_dirty_32 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  way0_dirty_33 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  way0_dirty_34 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  way0_dirty_35 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  way0_dirty_36 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  way0_dirty_37 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  way0_dirty_38 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  way0_dirty_39 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  way0_dirty_40 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  way0_dirty_41 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  way0_dirty_42 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  way0_dirty_43 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  way0_dirty_44 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  way0_dirty_45 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  way0_dirty_46 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  way0_dirty_47 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  way0_dirty_48 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  way0_dirty_49 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  way0_dirty_50 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  way0_dirty_51 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  way0_dirty_52 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  way0_dirty_53 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  way0_dirty_54 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  way0_dirty_55 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  way0_dirty_56 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  way0_dirty_57 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  way0_dirty_58 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  way0_dirty_59 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  way0_dirty_60 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  way0_dirty_61 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  way0_dirty_62 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  way0_dirty_63 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  way0_dirty_64 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  way0_dirty_65 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  way0_dirty_66 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  way0_dirty_67 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  way0_dirty_68 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  way0_dirty_69 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  way0_dirty_70 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  way0_dirty_71 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  way0_dirty_72 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  way0_dirty_73 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  way0_dirty_74 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  way0_dirty_75 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  way0_dirty_76 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  way0_dirty_77 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  way0_dirty_78 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  way0_dirty_79 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  way0_dirty_80 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  way0_dirty_81 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  way0_dirty_82 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  way0_dirty_83 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  way0_dirty_84 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  way0_dirty_85 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  way0_dirty_86 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  way0_dirty_87 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  way0_dirty_88 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  way0_dirty_89 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  way0_dirty_90 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  way0_dirty_91 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  way0_dirty_92 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  way0_dirty_93 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  way0_dirty_94 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  way0_dirty_95 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  way0_dirty_96 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  way0_dirty_97 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  way0_dirty_98 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  way0_dirty_99 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  way0_dirty_100 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  way0_dirty_101 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  way0_dirty_102 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  way0_dirty_103 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  way0_dirty_104 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  way0_dirty_105 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  way0_dirty_106 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  way0_dirty_107 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  way0_dirty_108 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  way0_dirty_109 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  way0_dirty_110 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  way0_dirty_111 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  way0_dirty_112 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  way0_dirty_113 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  way0_dirty_114 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  way0_dirty_115 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  way0_dirty_116 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  way0_dirty_117 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  way0_dirty_118 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  way0_dirty_119 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  way0_dirty_120 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  way0_dirty_121 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  way0_dirty_122 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  way0_dirty_123 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  way0_dirty_124 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  way0_dirty_125 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  way0_dirty_126 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  way0_dirty_127 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  way1_dirty_0 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  way1_dirty_1 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  way1_dirty_2 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  way1_dirty_3 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  way1_dirty_4 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  way1_dirty_5 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  way1_dirty_6 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  way1_dirty_7 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  way1_dirty_8 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  way1_dirty_9 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  way1_dirty_10 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  way1_dirty_11 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  way1_dirty_12 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  way1_dirty_13 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  way1_dirty_14 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  way1_dirty_15 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  way1_dirty_16 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  way1_dirty_17 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  way1_dirty_18 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  way1_dirty_19 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  way1_dirty_20 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  way1_dirty_21 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  way1_dirty_22 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  way1_dirty_23 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  way1_dirty_24 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  way1_dirty_25 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  way1_dirty_26 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  way1_dirty_27 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  way1_dirty_28 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  way1_dirty_29 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  way1_dirty_30 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  way1_dirty_31 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  way1_dirty_32 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  way1_dirty_33 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  way1_dirty_34 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  way1_dirty_35 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  way1_dirty_36 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  way1_dirty_37 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  way1_dirty_38 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  way1_dirty_39 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  way1_dirty_40 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  way1_dirty_41 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  way1_dirty_42 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  way1_dirty_43 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  way1_dirty_44 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  way1_dirty_45 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  way1_dirty_46 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  way1_dirty_47 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  way1_dirty_48 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  way1_dirty_49 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  way1_dirty_50 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  way1_dirty_51 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  way1_dirty_52 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  way1_dirty_53 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  way1_dirty_54 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  way1_dirty_55 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  way1_dirty_56 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  way1_dirty_57 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  way1_dirty_58 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  way1_dirty_59 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  way1_dirty_60 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  way1_dirty_61 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  way1_dirty_62 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  way1_dirty_63 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  way1_dirty_64 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  way1_dirty_65 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  way1_dirty_66 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  way1_dirty_67 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  way1_dirty_68 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  way1_dirty_69 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  way1_dirty_70 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  way1_dirty_71 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  way1_dirty_72 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  way1_dirty_73 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  way1_dirty_74 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  way1_dirty_75 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  way1_dirty_76 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  way1_dirty_77 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  way1_dirty_78 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  way1_dirty_79 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  way1_dirty_80 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  way1_dirty_81 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  way1_dirty_82 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  way1_dirty_83 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  way1_dirty_84 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  way1_dirty_85 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  way1_dirty_86 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  way1_dirty_87 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  way1_dirty_88 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  way1_dirty_89 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  way1_dirty_90 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  way1_dirty_91 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  way1_dirty_92 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  way1_dirty_93 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  way1_dirty_94 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  way1_dirty_95 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  way1_dirty_96 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  way1_dirty_97 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  way1_dirty_98 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  way1_dirty_99 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  way1_dirty_100 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  way1_dirty_101 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  way1_dirty_102 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  way1_dirty_103 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  way1_dirty_104 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  way1_dirty_105 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  way1_dirty_106 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  way1_dirty_107 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  way1_dirty_108 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  way1_dirty_109 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  way1_dirty_110 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  way1_dirty_111 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  way1_dirty_112 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  way1_dirty_113 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  way1_dirty_114 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  way1_dirty_115 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  way1_dirty_116 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  way1_dirty_117 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  way1_dirty_118 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  way1_dirty_119 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  way1_dirty_120 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  way1_dirty_121 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  way1_dirty_122 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  way1_dirty_123 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  way1_dirty_124 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  way1_dirty_125 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  way1_dirty_126 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  way1_dirty_127 = _RAND_387[0:0];
  _RAND_388 = {2{`RANDOM}};
  stage1_addr_line_mapping = _RAND_388[63:0];
  _RAND_389 = {1{`RANDOM}};
  stage1_sram_cache_reg = _RAND_389[0:0];
  _RAND_390 = {2{`RANDOM}};
  stage1_sram_wdata_reg = _RAND_390[63:0];
  _RAND_391 = {1{`RANDOM}};
  stage1_sram_size_reg = _RAND_391[1:0];
  _RAND_392 = {1{`RANDOM}};
  stage1_sram_wr_reg = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  stage1_sram_req_reg = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  stage1_sram_hit0_reg = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  stage1_sram_hit1_reg = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  stage1_sram_valid0_reg = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  stage1_sram_valid1_reg = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  stage1_wstrb_reg = _RAND_398[7:0];
  _RAND_399 = {2{`RANDOM}};
  stage1_sram_phy_addr_reg = _RAND_399[63:0];
  _RAND_400 = {1{`RANDOM}};
  data_write_back_counter = _RAND_400[7:0];
  _RAND_401 = {1{`RANDOM}};
  stage2_sram_write_reg = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  stage1_stall_reg = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  write_access_complete_reg = _RAND_403[0:0];
  _RAND_404 = {2{`RANDOM}};
  stage2_sram_addr_reg = _RAND_404[63:0];
  _RAND_405 = {1{`RANDOM}};
  stage2_hit0_reg = _RAND_405[0:0];
  _RAND_406 = {2{`RANDOM}};
  sram_rdata_reg = _RAND_406[63:0];
  _RAND_407 = {1{`RANDOM}};
  stage2_stall_reg = _RAND_407[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    work_state = 5'h18;
  end
  if (reset) begin
    write_counter = 3'h0;
  end
  if (reset) begin
    read_counter = 3'h0;
  end
  if (reset) begin
    wait_data = 64'h0;
  end
  if (reset) begin
    lru_0 = 1'h0;
  end
  if (reset) begin
    lru_1 = 1'h0;
  end
  if (reset) begin
    lru_2 = 1'h0;
  end
  if (reset) begin
    lru_3 = 1'h0;
  end
  if (reset) begin
    lru_4 = 1'h0;
  end
  if (reset) begin
    lru_5 = 1'h0;
  end
  if (reset) begin
    lru_6 = 1'h0;
  end
  if (reset) begin
    lru_7 = 1'h0;
  end
  if (reset) begin
    lru_8 = 1'h0;
  end
  if (reset) begin
    lru_9 = 1'h0;
  end
  if (reset) begin
    lru_10 = 1'h0;
  end
  if (reset) begin
    lru_11 = 1'h0;
  end
  if (reset) begin
    lru_12 = 1'h0;
  end
  if (reset) begin
    lru_13 = 1'h0;
  end
  if (reset) begin
    lru_14 = 1'h0;
  end
  if (reset) begin
    lru_15 = 1'h0;
  end
  if (reset) begin
    lru_16 = 1'h0;
  end
  if (reset) begin
    lru_17 = 1'h0;
  end
  if (reset) begin
    lru_18 = 1'h0;
  end
  if (reset) begin
    lru_19 = 1'h0;
  end
  if (reset) begin
    lru_20 = 1'h0;
  end
  if (reset) begin
    lru_21 = 1'h0;
  end
  if (reset) begin
    lru_22 = 1'h0;
  end
  if (reset) begin
    lru_23 = 1'h0;
  end
  if (reset) begin
    lru_24 = 1'h0;
  end
  if (reset) begin
    lru_25 = 1'h0;
  end
  if (reset) begin
    lru_26 = 1'h0;
  end
  if (reset) begin
    lru_27 = 1'h0;
  end
  if (reset) begin
    lru_28 = 1'h0;
  end
  if (reset) begin
    lru_29 = 1'h0;
  end
  if (reset) begin
    lru_30 = 1'h0;
  end
  if (reset) begin
    lru_31 = 1'h0;
  end
  if (reset) begin
    lru_32 = 1'h0;
  end
  if (reset) begin
    lru_33 = 1'h0;
  end
  if (reset) begin
    lru_34 = 1'h0;
  end
  if (reset) begin
    lru_35 = 1'h0;
  end
  if (reset) begin
    lru_36 = 1'h0;
  end
  if (reset) begin
    lru_37 = 1'h0;
  end
  if (reset) begin
    lru_38 = 1'h0;
  end
  if (reset) begin
    lru_39 = 1'h0;
  end
  if (reset) begin
    lru_40 = 1'h0;
  end
  if (reset) begin
    lru_41 = 1'h0;
  end
  if (reset) begin
    lru_42 = 1'h0;
  end
  if (reset) begin
    lru_43 = 1'h0;
  end
  if (reset) begin
    lru_44 = 1'h0;
  end
  if (reset) begin
    lru_45 = 1'h0;
  end
  if (reset) begin
    lru_46 = 1'h0;
  end
  if (reset) begin
    lru_47 = 1'h0;
  end
  if (reset) begin
    lru_48 = 1'h0;
  end
  if (reset) begin
    lru_49 = 1'h0;
  end
  if (reset) begin
    lru_50 = 1'h0;
  end
  if (reset) begin
    lru_51 = 1'h0;
  end
  if (reset) begin
    lru_52 = 1'h0;
  end
  if (reset) begin
    lru_53 = 1'h0;
  end
  if (reset) begin
    lru_54 = 1'h0;
  end
  if (reset) begin
    lru_55 = 1'h0;
  end
  if (reset) begin
    lru_56 = 1'h0;
  end
  if (reset) begin
    lru_57 = 1'h0;
  end
  if (reset) begin
    lru_58 = 1'h0;
  end
  if (reset) begin
    lru_59 = 1'h0;
  end
  if (reset) begin
    lru_60 = 1'h0;
  end
  if (reset) begin
    lru_61 = 1'h0;
  end
  if (reset) begin
    lru_62 = 1'h0;
  end
  if (reset) begin
    lru_63 = 1'h0;
  end
  if (reset) begin
    lru_64 = 1'h0;
  end
  if (reset) begin
    lru_65 = 1'h0;
  end
  if (reset) begin
    lru_66 = 1'h0;
  end
  if (reset) begin
    lru_67 = 1'h0;
  end
  if (reset) begin
    lru_68 = 1'h0;
  end
  if (reset) begin
    lru_69 = 1'h0;
  end
  if (reset) begin
    lru_70 = 1'h0;
  end
  if (reset) begin
    lru_71 = 1'h0;
  end
  if (reset) begin
    lru_72 = 1'h0;
  end
  if (reset) begin
    lru_73 = 1'h0;
  end
  if (reset) begin
    lru_74 = 1'h0;
  end
  if (reset) begin
    lru_75 = 1'h0;
  end
  if (reset) begin
    lru_76 = 1'h0;
  end
  if (reset) begin
    lru_77 = 1'h0;
  end
  if (reset) begin
    lru_78 = 1'h0;
  end
  if (reset) begin
    lru_79 = 1'h0;
  end
  if (reset) begin
    lru_80 = 1'h0;
  end
  if (reset) begin
    lru_81 = 1'h0;
  end
  if (reset) begin
    lru_82 = 1'h0;
  end
  if (reset) begin
    lru_83 = 1'h0;
  end
  if (reset) begin
    lru_84 = 1'h0;
  end
  if (reset) begin
    lru_85 = 1'h0;
  end
  if (reset) begin
    lru_86 = 1'h0;
  end
  if (reset) begin
    lru_87 = 1'h0;
  end
  if (reset) begin
    lru_88 = 1'h0;
  end
  if (reset) begin
    lru_89 = 1'h0;
  end
  if (reset) begin
    lru_90 = 1'h0;
  end
  if (reset) begin
    lru_91 = 1'h0;
  end
  if (reset) begin
    lru_92 = 1'h0;
  end
  if (reset) begin
    lru_93 = 1'h0;
  end
  if (reset) begin
    lru_94 = 1'h0;
  end
  if (reset) begin
    lru_95 = 1'h0;
  end
  if (reset) begin
    lru_96 = 1'h0;
  end
  if (reset) begin
    lru_97 = 1'h0;
  end
  if (reset) begin
    lru_98 = 1'h0;
  end
  if (reset) begin
    lru_99 = 1'h0;
  end
  if (reset) begin
    lru_100 = 1'h0;
  end
  if (reset) begin
    lru_101 = 1'h0;
  end
  if (reset) begin
    lru_102 = 1'h0;
  end
  if (reset) begin
    lru_103 = 1'h0;
  end
  if (reset) begin
    lru_104 = 1'h0;
  end
  if (reset) begin
    lru_105 = 1'h0;
  end
  if (reset) begin
    lru_106 = 1'h0;
  end
  if (reset) begin
    lru_107 = 1'h0;
  end
  if (reset) begin
    lru_108 = 1'h0;
  end
  if (reset) begin
    lru_109 = 1'h0;
  end
  if (reset) begin
    lru_110 = 1'h0;
  end
  if (reset) begin
    lru_111 = 1'h0;
  end
  if (reset) begin
    lru_112 = 1'h0;
  end
  if (reset) begin
    lru_113 = 1'h0;
  end
  if (reset) begin
    lru_114 = 1'h0;
  end
  if (reset) begin
    lru_115 = 1'h0;
  end
  if (reset) begin
    lru_116 = 1'h0;
  end
  if (reset) begin
    lru_117 = 1'h0;
  end
  if (reset) begin
    lru_118 = 1'h0;
  end
  if (reset) begin
    lru_119 = 1'h0;
  end
  if (reset) begin
    lru_120 = 1'h0;
  end
  if (reset) begin
    lru_121 = 1'h0;
  end
  if (reset) begin
    lru_122 = 1'h0;
  end
  if (reset) begin
    lru_123 = 1'h0;
  end
  if (reset) begin
    lru_124 = 1'h0;
  end
  if (reset) begin
    lru_125 = 1'h0;
  end
  if (reset) begin
    lru_126 = 1'h0;
  end
  if (reset) begin
    lru_127 = 1'h0;
  end
  if (reset) begin
    way0_dirty_0 = 1'h0;
  end
  if (reset) begin
    way0_dirty_1 = 1'h0;
  end
  if (reset) begin
    way0_dirty_2 = 1'h0;
  end
  if (reset) begin
    way0_dirty_3 = 1'h0;
  end
  if (reset) begin
    way0_dirty_4 = 1'h0;
  end
  if (reset) begin
    way0_dirty_5 = 1'h0;
  end
  if (reset) begin
    way0_dirty_6 = 1'h0;
  end
  if (reset) begin
    way0_dirty_7 = 1'h0;
  end
  if (reset) begin
    way0_dirty_8 = 1'h0;
  end
  if (reset) begin
    way0_dirty_9 = 1'h0;
  end
  if (reset) begin
    way0_dirty_10 = 1'h0;
  end
  if (reset) begin
    way0_dirty_11 = 1'h0;
  end
  if (reset) begin
    way0_dirty_12 = 1'h0;
  end
  if (reset) begin
    way0_dirty_13 = 1'h0;
  end
  if (reset) begin
    way0_dirty_14 = 1'h0;
  end
  if (reset) begin
    way0_dirty_15 = 1'h0;
  end
  if (reset) begin
    way0_dirty_16 = 1'h0;
  end
  if (reset) begin
    way0_dirty_17 = 1'h0;
  end
  if (reset) begin
    way0_dirty_18 = 1'h0;
  end
  if (reset) begin
    way0_dirty_19 = 1'h0;
  end
  if (reset) begin
    way0_dirty_20 = 1'h0;
  end
  if (reset) begin
    way0_dirty_21 = 1'h0;
  end
  if (reset) begin
    way0_dirty_22 = 1'h0;
  end
  if (reset) begin
    way0_dirty_23 = 1'h0;
  end
  if (reset) begin
    way0_dirty_24 = 1'h0;
  end
  if (reset) begin
    way0_dirty_25 = 1'h0;
  end
  if (reset) begin
    way0_dirty_26 = 1'h0;
  end
  if (reset) begin
    way0_dirty_27 = 1'h0;
  end
  if (reset) begin
    way0_dirty_28 = 1'h0;
  end
  if (reset) begin
    way0_dirty_29 = 1'h0;
  end
  if (reset) begin
    way0_dirty_30 = 1'h0;
  end
  if (reset) begin
    way0_dirty_31 = 1'h0;
  end
  if (reset) begin
    way0_dirty_32 = 1'h0;
  end
  if (reset) begin
    way0_dirty_33 = 1'h0;
  end
  if (reset) begin
    way0_dirty_34 = 1'h0;
  end
  if (reset) begin
    way0_dirty_35 = 1'h0;
  end
  if (reset) begin
    way0_dirty_36 = 1'h0;
  end
  if (reset) begin
    way0_dirty_37 = 1'h0;
  end
  if (reset) begin
    way0_dirty_38 = 1'h0;
  end
  if (reset) begin
    way0_dirty_39 = 1'h0;
  end
  if (reset) begin
    way0_dirty_40 = 1'h0;
  end
  if (reset) begin
    way0_dirty_41 = 1'h0;
  end
  if (reset) begin
    way0_dirty_42 = 1'h0;
  end
  if (reset) begin
    way0_dirty_43 = 1'h0;
  end
  if (reset) begin
    way0_dirty_44 = 1'h0;
  end
  if (reset) begin
    way0_dirty_45 = 1'h0;
  end
  if (reset) begin
    way0_dirty_46 = 1'h0;
  end
  if (reset) begin
    way0_dirty_47 = 1'h0;
  end
  if (reset) begin
    way0_dirty_48 = 1'h0;
  end
  if (reset) begin
    way0_dirty_49 = 1'h0;
  end
  if (reset) begin
    way0_dirty_50 = 1'h0;
  end
  if (reset) begin
    way0_dirty_51 = 1'h0;
  end
  if (reset) begin
    way0_dirty_52 = 1'h0;
  end
  if (reset) begin
    way0_dirty_53 = 1'h0;
  end
  if (reset) begin
    way0_dirty_54 = 1'h0;
  end
  if (reset) begin
    way0_dirty_55 = 1'h0;
  end
  if (reset) begin
    way0_dirty_56 = 1'h0;
  end
  if (reset) begin
    way0_dirty_57 = 1'h0;
  end
  if (reset) begin
    way0_dirty_58 = 1'h0;
  end
  if (reset) begin
    way0_dirty_59 = 1'h0;
  end
  if (reset) begin
    way0_dirty_60 = 1'h0;
  end
  if (reset) begin
    way0_dirty_61 = 1'h0;
  end
  if (reset) begin
    way0_dirty_62 = 1'h0;
  end
  if (reset) begin
    way0_dirty_63 = 1'h0;
  end
  if (reset) begin
    way0_dirty_64 = 1'h0;
  end
  if (reset) begin
    way0_dirty_65 = 1'h0;
  end
  if (reset) begin
    way0_dirty_66 = 1'h0;
  end
  if (reset) begin
    way0_dirty_67 = 1'h0;
  end
  if (reset) begin
    way0_dirty_68 = 1'h0;
  end
  if (reset) begin
    way0_dirty_69 = 1'h0;
  end
  if (reset) begin
    way0_dirty_70 = 1'h0;
  end
  if (reset) begin
    way0_dirty_71 = 1'h0;
  end
  if (reset) begin
    way0_dirty_72 = 1'h0;
  end
  if (reset) begin
    way0_dirty_73 = 1'h0;
  end
  if (reset) begin
    way0_dirty_74 = 1'h0;
  end
  if (reset) begin
    way0_dirty_75 = 1'h0;
  end
  if (reset) begin
    way0_dirty_76 = 1'h0;
  end
  if (reset) begin
    way0_dirty_77 = 1'h0;
  end
  if (reset) begin
    way0_dirty_78 = 1'h0;
  end
  if (reset) begin
    way0_dirty_79 = 1'h0;
  end
  if (reset) begin
    way0_dirty_80 = 1'h0;
  end
  if (reset) begin
    way0_dirty_81 = 1'h0;
  end
  if (reset) begin
    way0_dirty_82 = 1'h0;
  end
  if (reset) begin
    way0_dirty_83 = 1'h0;
  end
  if (reset) begin
    way0_dirty_84 = 1'h0;
  end
  if (reset) begin
    way0_dirty_85 = 1'h0;
  end
  if (reset) begin
    way0_dirty_86 = 1'h0;
  end
  if (reset) begin
    way0_dirty_87 = 1'h0;
  end
  if (reset) begin
    way0_dirty_88 = 1'h0;
  end
  if (reset) begin
    way0_dirty_89 = 1'h0;
  end
  if (reset) begin
    way0_dirty_90 = 1'h0;
  end
  if (reset) begin
    way0_dirty_91 = 1'h0;
  end
  if (reset) begin
    way0_dirty_92 = 1'h0;
  end
  if (reset) begin
    way0_dirty_93 = 1'h0;
  end
  if (reset) begin
    way0_dirty_94 = 1'h0;
  end
  if (reset) begin
    way0_dirty_95 = 1'h0;
  end
  if (reset) begin
    way0_dirty_96 = 1'h0;
  end
  if (reset) begin
    way0_dirty_97 = 1'h0;
  end
  if (reset) begin
    way0_dirty_98 = 1'h0;
  end
  if (reset) begin
    way0_dirty_99 = 1'h0;
  end
  if (reset) begin
    way0_dirty_100 = 1'h0;
  end
  if (reset) begin
    way0_dirty_101 = 1'h0;
  end
  if (reset) begin
    way0_dirty_102 = 1'h0;
  end
  if (reset) begin
    way0_dirty_103 = 1'h0;
  end
  if (reset) begin
    way0_dirty_104 = 1'h0;
  end
  if (reset) begin
    way0_dirty_105 = 1'h0;
  end
  if (reset) begin
    way0_dirty_106 = 1'h0;
  end
  if (reset) begin
    way0_dirty_107 = 1'h0;
  end
  if (reset) begin
    way0_dirty_108 = 1'h0;
  end
  if (reset) begin
    way0_dirty_109 = 1'h0;
  end
  if (reset) begin
    way0_dirty_110 = 1'h0;
  end
  if (reset) begin
    way0_dirty_111 = 1'h0;
  end
  if (reset) begin
    way0_dirty_112 = 1'h0;
  end
  if (reset) begin
    way0_dirty_113 = 1'h0;
  end
  if (reset) begin
    way0_dirty_114 = 1'h0;
  end
  if (reset) begin
    way0_dirty_115 = 1'h0;
  end
  if (reset) begin
    way0_dirty_116 = 1'h0;
  end
  if (reset) begin
    way0_dirty_117 = 1'h0;
  end
  if (reset) begin
    way0_dirty_118 = 1'h0;
  end
  if (reset) begin
    way0_dirty_119 = 1'h0;
  end
  if (reset) begin
    way0_dirty_120 = 1'h0;
  end
  if (reset) begin
    way0_dirty_121 = 1'h0;
  end
  if (reset) begin
    way0_dirty_122 = 1'h0;
  end
  if (reset) begin
    way0_dirty_123 = 1'h0;
  end
  if (reset) begin
    way0_dirty_124 = 1'h0;
  end
  if (reset) begin
    way0_dirty_125 = 1'h0;
  end
  if (reset) begin
    way0_dirty_126 = 1'h0;
  end
  if (reset) begin
    way0_dirty_127 = 1'h0;
  end
  if (reset) begin
    way1_dirty_0 = 1'h0;
  end
  if (reset) begin
    way1_dirty_1 = 1'h0;
  end
  if (reset) begin
    way1_dirty_2 = 1'h0;
  end
  if (reset) begin
    way1_dirty_3 = 1'h0;
  end
  if (reset) begin
    way1_dirty_4 = 1'h0;
  end
  if (reset) begin
    way1_dirty_5 = 1'h0;
  end
  if (reset) begin
    way1_dirty_6 = 1'h0;
  end
  if (reset) begin
    way1_dirty_7 = 1'h0;
  end
  if (reset) begin
    way1_dirty_8 = 1'h0;
  end
  if (reset) begin
    way1_dirty_9 = 1'h0;
  end
  if (reset) begin
    way1_dirty_10 = 1'h0;
  end
  if (reset) begin
    way1_dirty_11 = 1'h0;
  end
  if (reset) begin
    way1_dirty_12 = 1'h0;
  end
  if (reset) begin
    way1_dirty_13 = 1'h0;
  end
  if (reset) begin
    way1_dirty_14 = 1'h0;
  end
  if (reset) begin
    way1_dirty_15 = 1'h0;
  end
  if (reset) begin
    way1_dirty_16 = 1'h0;
  end
  if (reset) begin
    way1_dirty_17 = 1'h0;
  end
  if (reset) begin
    way1_dirty_18 = 1'h0;
  end
  if (reset) begin
    way1_dirty_19 = 1'h0;
  end
  if (reset) begin
    way1_dirty_20 = 1'h0;
  end
  if (reset) begin
    way1_dirty_21 = 1'h0;
  end
  if (reset) begin
    way1_dirty_22 = 1'h0;
  end
  if (reset) begin
    way1_dirty_23 = 1'h0;
  end
  if (reset) begin
    way1_dirty_24 = 1'h0;
  end
  if (reset) begin
    way1_dirty_25 = 1'h0;
  end
  if (reset) begin
    way1_dirty_26 = 1'h0;
  end
  if (reset) begin
    way1_dirty_27 = 1'h0;
  end
  if (reset) begin
    way1_dirty_28 = 1'h0;
  end
  if (reset) begin
    way1_dirty_29 = 1'h0;
  end
  if (reset) begin
    way1_dirty_30 = 1'h0;
  end
  if (reset) begin
    way1_dirty_31 = 1'h0;
  end
  if (reset) begin
    way1_dirty_32 = 1'h0;
  end
  if (reset) begin
    way1_dirty_33 = 1'h0;
  end
  if (reset) begin
    way1_dirty_34 = 1'h0;
  end
  if (reset) begin
    way1_dirty_35 = 1'h0;
  end
  if (reset) begin
    way1_dirty_36 = 1'h0;
  end
  if (reset) begin
    way1_dirty_37 = 1'h0;
  end
  if (reset) begin
    way1_dirty_38 = 1'h0;
  end
  if (reset) begin
    way1_dirty_39 = 1'h0;
  end
  if (reset) begin
    way1_dirty_40 = 1'h0;
  end
  if (reset) begin
    way1_dirty_41 = 1'h0;
  end
  if (reset) begin
    way1_dirty_42 = 1'h0;
  end
  if (reset) begin
    way1_dirty_43 = 1'h0;
  end
  if (reset) begin
    way1_dirty_44 = 1'h0;
  end
  if (reset) begin
    way1_dirty_45 = 1'h0;
  end
  if (reset) begin
    way1_dirty_46 = 1'h0;
  end
  if (reset) begin
    way1_dirty_47 = 1'h0;
  end
  if (reset) begin
    way1_dirty_48 = 1'h0;
  end
  if (reset) begin
    way1_dirty_49 = 1'h0;
  end
  if (reset) begin
    way1_dirty_50 = 1'h0;
  end
  if (reset) begin
    way1_dirty_51 = 1'h0;
  end
  if (reset) begin
    way1_dirty_52 = 1'h0;
  end
  if (reset) begin
    way1_dirty_53 = 1'h0;
  end
  if (reset) begin
    way1_dirty_54 = 1'h0;
  end
  if (reset) begin
    way1_dirty_55 = 1'h0;
  end
  if (reset) begin
    way1_dirty_56 = 1'h0;
  end
  if (reset) begin
    way1_dirty_57 = 1'h0;
  end
  if (reset) begin
    way1_dirty_58 = 1'h0;
  end
  if (reset) begin
    way1_dirty_59 = 1'h0;
  end
  if (reset) begin
    way1_dirty_60 = 1'h0;
  end
  if (reset) begin
    way1_dirty_61 = 1'h0;
  end
  if (reset) begin
    way1_dirty_62 = 1'h0;
  end
  if (reset) begin
    way1_dirty_63 = 1'h0;
  end
  if (reset) begin
    way1_dirty_64 = 1'h0;
  end
  if (reset) begin
    way1_dirty_65 = 1'h0;
  end
  if (reset) begin
    way1_dirty_66 = 1'h0;
  end
  if (reset) begin
    way1_dirty_67 = 1'h0;
  end
  if (reset) begin
    way1_dirty_68 = 1'h0;
  end
  if (reset) begin
    way1_dirty_69 = 1'h0;
  end
  if (reset) begin
    way1_dirty_70 = 1'h0;
  end
  if (reset) begin
    way1_dirty_71 = 1'h0;
  end
  if (reset) begin
    way1_dirty_72 = 1'h0;
  end
  if (reset) begin
    way1_dirty_73 = 1'h0;
  end
  if (reset) begin
    way1_dirty_74 = 1'h0;
  end
  if (reset) begin
    way1_dirty_75 = 1'h0;
  end
  if (reset) begin
    way1_dirty_76 = 1'h0;
  end
  if (reset) begin
    way1_dirty_77 = 1'h0;
  end
  if (reset) begin
    way1_dirty_78 = 1'h0;
  end
  if (reset) begin
    way1_dirty_79 = 1'h0;
  end
  if (reset) begin
    way1_dirty_80 = 1'h0;
  end
  if (reset) begin
    way1_dirty_81 = 1'h0;
  end
  if (reset) begin
    way1_dirty_82 = 1'h0;
  end
  if (reset) begin
    way1_dirty_83 = 1'h0;
  end
  if (reset) begin
    way1_dirty_84 = 1'h0;
  end
  if (reset) begin
    way1_dirty_85 = 1'h0;
  end
  if (reset) begin
    way1_dirty_86 = 1'h0;
  end
  if (reset) begin
    way1_dirty_87 = 1'h0;
  end
  if (reset) begin
    way1_dirty_88 = 1'h0;
  end
  if (reset) begin
    way1_dirty_89 = 1'h0;
  end
  if (reset) begin
    way1_dirty_90 = 1'h0;
  end
  if (reset) begin
    way1_dirty_91 = 1'h0;
  end
  if (reset) begin
    way1_dirty_92 = 1'h0;
  end
  if (reset) begin
    way1_dirty_93 = 1'h0;
  end
  if (reset) begin
    way1_dirty_94 = 1'h0;
  end
  if (reset) begin
    way1_dirty_95 = 1'h0;
  end
  if (reset) begin
    way1_dirty_96 = 1'h0;
  end
  if (reset) begin
    way1_dirty_97 = 1'h0;
  end
  if (reset) begin
    way1_dirty_98 = 1'h0;
  end
  if (reset) begin
    way1_dirty_99 = 1'h0;
  end
  if (reset) begin
    way1_dirty_100 = 1'h0;
  end
  if (reset) begin
    way1_dirty_101 = 1'h0;
  end
  if (reset) begin
    way1_dirty_102 = 1'h0;
  end
  if (reset) begin
    way1_dirty_103 = 1'h0;
  end
  if (reset) begin
    way1_dirty_104 = 1'h0;
  end
  if (reset) begin
    way1_dirty_105 = 1'h0;
  end
  if (reset) begin
    way1_dirty_106 = 1'h0;
  end
  if (reset) begin
    way1_dirty_107 = 1'h0;
  end
  if (reset) begin
    way1_dirty_108 = 1'h0;
  end
  if (reset) begin
    way1_dirty_109 = 1'h0;
  end
  if (reset) begin
    way1_dirty_110 = 1'h0;
  end
  if (reset) begin
    way1_dirty_111 = 1'h0;
  end
  if (reset) begin
    way1_dirty_112 = 1'h0;
  end
  if (reset) begin
    way1_dirty_113 = 1'h0;
  end
  if (reset) begin
    way1_dirty_114 = 1'h0;
  end
  if (reset) begin
    way1_dirty_115 = 1'h0;
  end
  if (reset) begin
    way1_dirty_116 = 1'h0;
  end
  if (reset) begin
    way1_dirty_117 = 1'h0;
  end
  if (reset) begin
    way1_dirty_118 = 1'h0;
  end
  if (reset) begin
    way1_dirty_119 = 1'h0;
  end
  if (reset) begin
    way1_dirty_120 = 1'h0;
  end
  if (reset) begin
    way1_dirty_121 = 1'h0;
  end
  if (reset) begin
    way1_dirty_122 = 1'h0;
  end
  if (reset) begin
    way1_dirty_123 = 1'h0;
  end
  if (reset) begin
    way1_dirty_124 = 1'h0;
  end
  if (reset) begin
    way1_dirty_125 = 1'h0;
  end
  if (reset) begin
    way1_dirty_126 = 1'h0;
  end
  if (reset) begin
    way1_dirty_127 = 1'h0;
  end
  if (reset) begin
    stage1_addr_line_mapping = 64'h0;
  end
  if (reset) begin
    stage1_sram_cache_reg = 1'h0;
  end
  if (reset) begin
    stage1_sram_wdata_reg = 64'h0;
  end
  if (reset) begin
    stage1_sram_size_reg = 2'h0;
  end
  if (reset) begin
    stage1_sram_wr_reg = 1'h0;
  end
  if (reset) begin
    stage1_sram_req_reg = 1'h0;
  end
  if (reset) begin
    stage1_sram_hit0_reg = 1'h0;
  end
  if (reset) begin
    stage1_sram_hit1_reg = 1'h0;
  end
  if (reset) begin
    stage1_sram_valid0_reg = 1'h0;
  end
  if (reset) begin
    stage1_sram_valid1_reg = 1'h0;
  end
  if (reset) begin
    stage1_wstrb_reg = 8'h0;
  end
  if (reset) begin
    stage1_sram_phy_addr_reg = 64'h0;
  end
  if (reset) begin
    data_write_back_counter = 8'h0;
  end
  if (reset) begin
    stage2_sram_write_reg = 1'h0;
  end
  if (reset) begin
    stage1_stall_reg = 1'h0;
  end
  if (reset) begin
    write_access_complete_reg = 1'h0;
  end
  if (reset) begin
    stage2_sram_addr_reg = 64'h0;
  end
  if (reset) begin
    stage2_hit0_reg = 1'h0;
  end
  if (reset) begin
    sram_rdata_reg = 64'h0;
  end
  if (reset) begin
    stage2_stall_reg = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module axi_cross_bar(
  input         clock,
  input         reset,
  input  [63:0] io_m_port_0_araddr,
  input  [3:0]  io_m_port_0_arlen,
  input  [1:0]  io_m_port_0_arburst,
  input         io_m_port_0_arvalid,
  output        io_m_port_0_arready,
  output [63:0] io_m_port_0_rdata,
  output        io_m_port_0_rlast,
  output        io_m_port_0_rvalid,
  input  [63:0] io_m_port_1_araddr,
  input  [3:0]  io_m_port_1_arlen,
  input  [2:0]  io_m_port_1_arsize,
  input  [1:0]  io_m_port_1_arburst,
  input         io_m_port_1_arvalid,
  output        io_m_port_1_arready,
  output [63:0] io_m_port_1_rdata,
  output        io_m_port_1_rlast,
  output        io_m_port_1_rvalid,
  input  [63:0] io_m_port_1_awaddr,
  input  [3:0]  io_m_port_1_awlen,
  input  [2:0]  io_m_port_1_awsize,
  input  [1:0]  io_m_port_1_awburst,
  input         io_m_port_1_awvalid,
  output        io_m_port_1_awready,
  input  [63:0] io_m_port_1_wdata,
  input  [7:0]  io_m_port_1_wstrb,
  input         io_m_port_1_wlast,
  input         io_m_port_1_wvalid,
  output        io_m_port_1_wready,
  output        io_m_port_1_bvalid,
  output [3:0]  io_s_port_arid,
  output [63:0] io_s_port_araddr,
  output [3:0]  io_s_port_arlen,
  output [2:0]  io_s_port_arsize,
  output [1:0]  io_s_port_arburst,
  output        io_s_port_arvalid,
  input         io_s_port_arready,
  input  [63:0] io_s_port_rdata,
  input         io_s_port_rlast,
  input         io_s_port_rvalid,
  output        io_s_port_rready,
  output [3:0]  io_s_port_awid,
  output [63:0] io_s_port_awaddr,
  output [3:0]  io_s_port_awlen,
  output [2:0]  io_s_port_awsize,
  output [1:0]  io_s_port_awburst,
  output        io_s_port_awvalid,
  input         io_s_port_awready,
  output [3:0]  io_s_port_wid,
  output [63:0] io_s_port_wdata,
  output [7:0]  io_s_port_wstrb,
  output        io_s_port_wlast,
  output        io_s_port_wvalid,
  input         io_s_port_wready,
  input         io_s_port_bvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg  r_inuse_0; // @[axi_ram_port.scala 119:30]
  reg  r_inuse_1; // @[axi_ram_port.scala 119:30]
  reg  w_inuse_1; // @[axi_ram_port.scala 121:30]
  wire [1:0] _T_3 = {w_inuse_1,1'h0}; // @[axi_ram_port.scala 125:93]
  wire  _GEN_4 = io_s_port_bvalid & w_inuse_1 ? 1'h0 : w_inuse_1; // @[axi_ram_port.scala 128:67 129:41 131:41]
  wire  w_inuse_wire_1 = (io_m_port_1_awvalid | io_m_port_1_wvalid) & _T_3 == 2'h0 | _GEN_4; // @[axi_ram_port.scala 125:110 127:41]
  wire [1:0] _w_inuse_0_T = {w_inuse_wire_1,1'h0}; // @[axi_ram_port.scala 139:48]
  wire [1:0] _w_inuse_0_T_6 = 2'h2 - 2'h1; // @[axi_ram_port.scala 139:117]
  wire  _w_inuse_0_T_7 = 2'h0 == _w_inuse_0_T_6; // @[axi_ram_port.scala 139:95]
  wire [1:0] _T_11 = {r_inuse_1,r_inuse_0}; // @[axi_ram_port.scala 141:93]
  wire  _GEN_2 = io_s_port_rlast & r_inuse_0 ? 1'h0 : r_inuse_0; // @[axi_ram_port.scala 143:65 144:41 146:41]
  wire  r_inuse_wire_0 = (io_m_port_0_arvalid | io_m_port_0_rvalid) & _T_11 == 2'h0 | _GEN_2; // @[axi_ram_port.scala 141:110 142:41]
  wire  _GEN_6 = io_s_port_rlast & r_inuse_1 ? 1'h0 : r_inuse_1; // @[axi_ram_port.scala 143:65 144:41 146:41]
  wire  r_inuse_wire_1 = (io_m_port_1_arvalid | io_m_port_1_rvalid) & _T_11 == 2'h0 | _GEN_6; // @[axi_ram_port.scala 141:110 142:41]
  wire [1:0] _r_inuse_0_T = {r_inuse_wire_1,r_inuse_wire_0}; // @[axi_ram_port.scala 156:49]
  wire [1:0] _r_inuse_0_T_3 = {{1'd0}, _r_inuse_0_T[1]}; // @[axi_ram_port.scala 156:56]
  wire  _w_inuse_1_T_7 = 2'h1 == _w_inuse_0_T_6; // @[axi_ram_port.scala 139:95]
  wire [1:0] _r_select_port_T_93 = r_inuse_0 ? io_m_port_0_arburst : 2'h0; // @[Mux.scala 27:73]
  wire [1:0] _r_select_port_T_94 = r_inuse_1 ? io_m_port_1_arburst : 2'h0; // @[Mux.scala 27:73]
  wire [2:0] _r_select_port_T_96 = r_inuse_0 ? 3'h3 : 3'h0; // @[Mux.scala 27:73]
  wire [2:0] _r_select_port_T_97 = r_inuse_1 ? io_m_port_1_arsize : 3'h0; // @[Mux.scala 27:73]
  wire [3:0] _r_select_port_T_99 = r_inuse_0 ? io_m_port_0_arlen : 4'h0; // @[Mux.scala 27:73]
  wire [3:0] _r_select_port_T_100 = r_inuse_1 ? io_m_port_1_arlen : 4'h0; // @[Mux.scala 27:73]
  wire [63:0] _r_select_port_T_102 = r_inuse_0 ? io_m_port_0_araddr : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _r_select_port_T_103 = r_inuse_1 ? io_m_port_1_araddr : 64'h0; // @[Mux.scala 27:73]
  assign io_m_port_0_arready = r_inuse_0 & io_s_port_arready; // @[axi_ram_port.scala 150:44]
  assign io_m_port_0_rdata = r_inuse_0 ? io_s_port_rdata : 64'h0; // @[axi_ram_port.scala 152:44]
  assign io_m_port_0_rlast = r_inuse_0 & io_s_port_rlast; // @[axi_ram_port.scala 154:44]
  assign io_m_port_0_rvalid = r_inuse_0 & io_s_port_rvalid; // @[axi_ram_port.scala 155:44]
  assign io_m_port_1_arready = r_inuse_1 & io_s_port_arready; // @[axi_ram_port.scala 150:44]
  assign io_m_port_1_rdata = r_inuse_1 ? io_s_port_rdata : 64'h0; // @[axi_ram_port.scala 152:44]
  assign io_m_port_1_rlast = r_inuse_1 & io_s_port_rlast; // @[axi_ram_port.scala 154:44]
  assign io_m_port_1_rvalid = r_inuse_1 & io_s_port_rvalid; // @[axi_ram_port.scala 155:44]
  assign io_m_port_1_awready = w_inuse_1 & io_s_port_awready; // @[axi_ram_port.scala 134:45]
  assign io_m_port_1_wready = w_inuse_1 & io_s_port_wready; // @[axi_ram_port.scala 135:45]
  assign io_m_port_1_bvalid = w_inuse_1 & io_s_port_bvalid; // @[axi_ram_port.scala 138:45]
  assign io_s_port_arid = r_inuse_1 ? 4'h1 : 4'h0; // @[Mux.scala 27:73]
  assign io_s_port_araddr = _r_select_port_T_102 | _r_select_port_T_103; // @[Mux.scala 27:73]
  assign io_s_port_arlen = _r_select_port_T_99 | _r_select_port_T_100; // @[Mux.scala 27:73]
  assign io_s_port_arsize = _r_select_port_T_96 | _r_select_port_T_97; // @[Mux.scala 27:73]
  assign io_s_port_arburst = _r_select_port_T_93 | _r_select_port_T_94; // @[Mux.scala 27:73]
  assign io_s_port_arvalid = r_inuse_0 & io_m_port_0_arvalid | r_inuse_1 & io_m_port_1_arvalid; // @[Mux.scala 27:73]
  assign io_s_port_rready = r_inuse_0 | r_inuse_1; // @[Mux.scala 27:73]
  assign io_s_port_awid = w_inuse_1 ? 4'h1 : 4'h0; // @[Mux.scala 27:73]
  assign io_s_port_awaddr = w_inuse_1 ? io_m_port_1_awaddr : 64'h0; // @[Mux.scala 27:73]
  assign io_s_port_awlen = w_inuse_1 ? io_m_port_1_awlen : 4'h0; // @[Mux.scala 27:73]
  assign io_s_port_awsize = w_inuse_1 ? io_m_port_1_awsize : 3'h0; // @[Mux.scala 27:73]
  assign io_s_port_awburst = w_inuse_1 ? io_m_port_1_awburst : 2'h0; // @[Mux.scala 27:73]
  assign io_s_port_awvalid = w_inuse_1 & io_m_port_1_awvalid; // @[Mux.scala 27:73]
  assign io_s_port_wid = w_inuse_1 ? 4'h1 : 4'h0; // @[Mux.scala 27:73]
  assign io_s_port_wdata = w_inuse_1 ? io_m_port_1_wdata : 64'h0; // @[Mux.scala 27:73]
  assign io_s_port_wstrb = w_inuse_1 ? io_m_port_1_wstrb : 8'h0; // @[Mux.scala 27:73]
  assign io_s_port_wlast = w_inuse_1 & io_m_port_1_wlast; // @[Mux.scala 27:73]
  assign io_s_port_wvalid = w_inuse_1 & io_m_port_1_wvalid; // @[Mux.scala 27:73]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[axi_ram_port.scala 156:34]
      r_inuse_0 <= 1'h0;
    end else begin
      r_inuse_0 <= (_r_inuse_0_T_3 == 2'h0 | _w_inuse_0_T_7) & r_inuse_wire_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[axi_ram_port.scala 156:34]
      r_inuse_1 <= 1'h0;
    end else begin
      r_inuse_1 <= (_r_inuse_0_T == 2'h0 | _w_inuse_1_T_7) & r_inuse_wire_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[axi_ram_port.scala 139:34]
      w_inuse_1 <= 1'h0;
    end else begin
      w_inuse_1 <= (_w_inuse_0_T == 2'h0 | 2'h1 == _w_inuse_0_T_6) & w_inuse_wire_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_inuse_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  r_inuse_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  w_inuse_1 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    r_inuse_0 = 1'h0;
  end
  if (reset) begin
    r_inuse_1 = 1'h0;
  end
  if (reset) begin
    w_inuse_1 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module axi_cross_bar_addr_switch(
  input         clock,
  input         reset,
  input  [63:0] io_m_port_0_araddr,
  input  [3:0]  io_m_port_0_arlen,
  input  [1:0]  io_m_port_0_arburst,
  input         io_m_port_0_arvalid,
  output        io_m_port_0_arready,
  output [63:0] io_m_port_0_rdata,
  output        io_m_port_0_rlast,
  output        io_m_port_0_rvalid,
  input  [63:0] io_m_port_1_araddr,
  input  [3:0]  io_m_port_1_arlen,
  input  [2:0]  io_m_port_1_arsize,
  input  [1:0]  io_m_port_1_arburst,
  input         io_m_port_1_arvalid,
  output        io_m_port_1_arready,
  output [63:0] io_m_port_1_rdata,
  output        io_m_port_1_rlast,
  output        io_m_port_1_rvalid,
  input  [63:0] io_m_port_1_awaddr,
  input  [3:0]  io_m_port_1_awlen,
  input  [2:0]  io_m_port_1_awsize,
  input  [1:0]  io_m_port_1_awburst,
  input         io_m_port_1_awvalid,
  output        io_m_port_1_awready,
  input  [63:0] io_m_port_1_wdata,
  input  [7:0]  io_m_port_1_wstrb,
  input         io_m_port_1_wlast,
  input         io_m_port_1_wvalid,
  output        io_m_port_1_wready,
  output        io_m_port_1_bvalid,
  output [3:0]  io_s_port_0_arid,
  output [63:0] io_s_port_0_araddr,
  output [3:0]  io_s_port_0_arlen,
  output [2:0]  io_s_port_0_arsize,
  output [1:0]  io_s_port_0_arburst,
  output        io_s_port_0_arvalid,
  input         io_s_port_0_arready,
  input  [63:0] io_s_port_0_rdata,
  input         io_s_port_0_rlast,
  input         io_s_port_0_rvalid,
  output        io_s_port_0_rready,
  output [3:0]  io_s_port_0_awid,
  output [63:0] io_s_port_0_awaddr,
  output [3:0]  io_s_port_0_awlen,
  output [2:0]  io_s_port_0_awsize,
  output [1:0]  io_s_port_0_awburst,
  output        io_s_port_0_awvalid,
  input         io_s_port_0_awready,
  output [3:0]  io_s_port_0_wid,
  output [63:0] io_s_port_0_wdata,
  output [7:0]  io_s_port_0_wstrb,
  output        io_s_port_0_wlast,
  output        io_s_port_0_wvalid,
  input         io_s_port_0_wready,
  input         io_s_port_0_bvalid,
  output        io_s_port_0_bready,
  output [63:0] io_s_port_1_araddr,
  output        io_s_port_1_arvalid,
  input  [63:0] io_s_port_1_rdata,
  input         io_s_port_1_rlast,
  input         io_s_port_1_rvalid,
  output        io_s_port_1_rready,
  output [63:0] io_s_port_1_awaddr,
  output [2:0]  io_s_port_1_awsize,
  output        io_s_port_1_awvalid,
  output [63:0] io_s_port_1_wdata,
  output        io_s_port_1_wvalid,
  input         io_s_port_1_wready,
  input         io_s_port_1_bvalid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  axi_cross_bar_clock; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_reset; // @[axi_ram_port.scala 204:38]
  wire [63:0] axi_cross_bar_io_m_port_0_araddr; // @[axi_ram_port.scala 204:38]
  wire [3:0] axi_cross_bar_io_m_port_0_arlen; // @[axi_ram_port.scala 204:38]
  wire [1:0] axi_cross_bar_io_m_port_0_arburst; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_m_port_0_arvalid; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_m_port_0_arready; // @[axi_ram_port.scala 204:38]
  wire [63:0] axi_cross_bar_io_m_port_0_rdata; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_m_port_0_rlast; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_m_port_0_rvalid; // @[axi_ram_port.scala 204:38]
  wire [63:0] axi_cross_bar_io_m_port_1_araddr; // @[axi_ram_port.scala 204:38]
  wire [3:0] axi_cross_bar_io_m_port_1_arlen; // @[axi_ram_port.scala 204:38]
  wire [2:0] axi_cross_bar_io_m_port_1_arsize; // @[axi_ram_port.scala 204:38]
  wire [1:0] axi_cross_bar_io_m_port_1_arburst; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_m_port_1_arvalid; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_m_port_1_arready; // @[axi_ram_port.scala 204:38]
  wire [63:0] axi_cross_bar_io_m_port_1_rdata; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_m_port_1_rlast; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_m_port_1_rvalid; // @[axi_ram_port.scala 204:38]
  wire [63:0] axi_cross_bar_io_m_port_1_awaddr; // @[axi_ram_port.scala 204:38]
  wire [3:0] axi_cross_bar_io_m_port_1_awlen; // @[axi_ram_port.scala 204:38]
  wire [2:0] axi_cross_bar_io_m_port_1_awsize; // @[axi_ram_port.scala 204:38]
  wire [1:0] axi_cross_bar_io_m_port_1_awburst; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_m_port_1_awvalid; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_m_port_1_awready; // @[axi_ram_port.scala 204:38]
  wire [63:0] axi_cross_bar_io_m_port_1_wdata; // @[axi_ram_port.scala 204:38]
  wire [7:0] axi_cross_bar_io_m_port_1_wstrb; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_m_port_1_wlast; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_m_port_1_wvalid; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_m_port_1_wready; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_m_port_1_bvalid; // @[axi_ram_port.scala 204:38]
  wire [3:0] axi_cross_bar_io_s_port_arid; // @[axi_ram_port.scala 204:38]
  wire [63:0] axi_cross_bar_io_s_port_araddr; // @[axi_ram_port.scala 204:38]
  wire [3:0] axi_cross_bar_io_s_port_arlen; // @[axi_ram_port.scala 204:38]
  wire [2:0] axi_cross_bar_io_s_port_arsize; // @[axi_ram_port.scala 204:38]
  wire [1:0] axi_cross_bar_io_s_port_arburst; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_s_port_arvalid; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_s_port_arready; // @[axi_ram_port.scala 204:38]
  wire [63:0] axi_cross_bar_io_s_port_rdata; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_s_port_rlast; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_s_port_rvalid; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_s_port_rready; // @[axi_ram_port.scala 204:38]
  wire [3:0] axi_cross_bar_io_s_port_awid; // @[axi_ram_port.scala 204:38]
  wire [63:0] axi_cross_bar_io_s_port_awaddr; // @[axi_ram_port.scala 204:38]
  wire [3:0] axi_cross_bar_io_s_port_awlen; // @[axi_ram_port.scala 204:38]
  wire [2:0] axi_cross_bar_io_s_port_awsize; // @[axi_ram_port.scala 204:38]
  wire [1:0] axi_cross_bar_io_s_port_awburst; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_s_port_awvalid; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_s_port_awready; // @[axi_ram_port.scala 204:38]
  wire [3:0] axi_cross_bar_io_s_port_wid; // @[axi_ram_port.scala 204:38]
  wire [63:0] axi_cross_bar_io_s_port_wdata; // @[axi_ram_port.scala 204:38]
  wire [7:0] axi_cross_bar_io_s_port_wstrb; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_s_port_wlast; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_s_port_wvalid; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_s_port_wready; // @[axi_ram_port.scala 204:38]
  wire  axi_cross_bar_io_s_port_bvalid; // @[axi_ram_port.scala 204:38]
  reg  select_s_port_num_r_0; // @[axi_ram_port.scala 209:43]
  reg  select_s_port_num_r_1; // @[axi_ram_port.scala 209:43]
  reg  select_s_port_num_w_0; // @[axi_ram_port.scala 210:43]
  reg  select_s_port_num_w_1; // @[axi_ram_port.scala 210:43]
  wire  _access_select_s_port_num_r_1_T = axi_cross_bar_io_s_port_arvalid; // @[axi_ram_port.scala 237:98]
  wire  _access_select_s_port_num_r_1_T_2 = axi_cross_bar_io_s_port_araddr < 64'h2000bfff; // @[axi_ram_port.scala 238:64]
  wire  _access_select_s_port_num_r_1_T_3 = axi_cross_bar_io_s_port_araddr >= 64'h20000000 &
    _access_select_s_port_num_r_1_T_2; // @[axi_ram_port.scala 237:182]
  wire  access_select_s_port_num_r_1 = axi_cross_bar_io_s_port_arvalid ? axi_cross_bar_io_s_port_araddr >= 64'h20000000
     & _access_select_s_port_num_r_1_T_2 : select_s_port_num_r_1; // @[axi_ram_port.scala 237:65]
  wire  _access_select_s_port_num_r_0_T_1 = ~access_select_s_port_num_r_1; // @[axi_ram_port.scala 219:90]
  wire  access_select_s_port_num_r_0 = _access_select_s_port_num_r_1_T ? _access_select_s_port_num_r_0_T_1 :
    select_s_port_num_r_0; // @[axi_ram_port.scala 218:69]
  wire [1:0] _r_to_be_T = {access_select_s_port_num_r_1,access_select_s_port_num_r_0}; // @[axi_ram_port.scala 217:78]
  wire  _access_select_s_port_num_w_1_T = axi_cross_bar_io_s_port_awvalid; // @[axi_ram_port.scala 242:98]
  wire  _access_select_s_port_num_w_1_T_2 = axi_cross_bar_io_s_port_awaddr < 64'h2000bfff; // @[axi_ram_port.scala 243:64]
  wire  _access_select_s_port_num_w_1_T_3 = axi_cross_bar_io_s_port_awaddr >= 64'h20000000 &
    _access_select_s_port_num_w_1_T_2; // @[axi_ram_port.scala 242:180]
  wire  access_select_s_port_num_w_1 = axi_cross_bar_io_s_port_awvalid ? axi_cross_bar_io_s_port_awaddr >= 64'h20000000
     & _access_select_s_port_num_w_1_T_2 : select_s_port_num_w_1; // @[axi_ram_port.scala 242:65]
  wire  _access_select_s_port_num_w_0_T_1 = ~access_select_s_port_num_w_1; // @[axi_ram_port.scala 223:90]
  wire  access_select_s_port_num_w_0 = _access_select_s_port_num_w_1_T ? _access_select_s_port_num_w_0_T_1 :
    select_s_port_num_w_0; // @[axi_ram_port.scala 222:73]
  wire [1:0] _w_to_be_T = {access_select_s_port_num_w_1,access_select_s_port_num_w_0}; // @[axi_ram_port.scala 221:78]
  wire [63:0] master_bundle_arready_0 = {{63'd0}, io_s_port_0_arready}; // @[axi_ram_port.scala 250:41 276:48]
  wire [63:0] _T_15 = access_select_s_port_num_r_0 ? master_bundle_arready_0 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_16 = access_select_s_port_num_r_1 ? 64'h1 : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_17 = _T_15 | _T_16; // @[Mux.scala 27:73]
  wire [63:0] _T_21 = access_select_s_port_num_r_0 ? io_s_port_0_rdata : 64'h0; // @[Mux.scala 27:73]
  wire [63:0] _T_22 = access_select_s_port_num_r_1 ? io_s_port_1_rdata : 64'h0; // @[Mux.scala 27:73]
  axi_cross_bar axi_cross_bar ( // @[axi_ram_port.scala 204:38]
    .clock(axi_cross_bar_clock),
    .reset(axi_cross_bar_reset),
    .io_m_port_0_araddr(axi_cross_bar_io_m_port_0_araddr),
    .io_m_port_0_arlen(axi_cross_bar_io_m_port_0_arlen),
    .io_m_port_0_arburst(axi_cross_bar_io_m_port_0_arburst),
    .io_m_port_0_arvalid(axi_cross_bar_io_m_port_0_arvalid),
    .io_m_port_0_arready(axi_cross_bar_io_m_port_0_arready),
    .io_m_port_0_rdata(axi_cross_bar_io_m_port_0_rdata),
    .io_m_port_0_rlast(axi_cross_bar_io_m_port_0_rlast),
    .io_m_port_0_rvalid(axi_cross_bar_io_m_port_0_rvalid),
    .io_m_port_1_araddr(axi_cross_bar_io_m_port_1_araddr),
    .io_m_port_1_arlen(axi_cross_bar_io_m_port_1_arlen),
    .io_m_port_1_arsize(axi_cross_bar_io_m_port_1_arsize),
    .io_m_port_1_arburst(axi_cross_bar_io_m_port_1_arburst),
    .io_m_port_1_arvalid(axi_cross_bar_io_m_port_1_arvalid),
    .io_m_port_1_arready(axi_cross_bar_io_m_port_1_arready),
    .io_m_port_1_rdata(axi_cross_bar_io_m_port_1_rdata),
    .io_m_port_1_rlast(axi_cross_bar_io_m_port_1_rlast),
    .io_m_port_1_rvalid(axi_cross_bar_io_m_port_1_rvalid),
    .io_m_port_1_awaddr(axi_cross_bar_io_m_port_1_awaddr),
    .io_m_port_1_awlen(axi_cross_bar_io_m_port_1_awlen),
    .io_m_port_1_awsize(axi_cross_bar_io_m_port_1_awsize),
    .io_m_port_1_awburst(axi_cross_bar_io_m_port_1_awburst),
    .io_m_port_1_awvalid(axi_cross_bar_io_m_port_1_awvalid),
    .io_m_port_1_awready(axi_cross_bar_io_m_port_1_awready),
    .io_m_port_1_wdata(axi_cross_bar_io_m_port_1_wdata),
    .io_m_port_1_wstrb(axi_cross_bar_io_m_port_1_wstrb),
    .io_m_port_1_wlast(axi_cross_bar_io_m_port_1_wlast),
    .io_m_port_1_wvalid(axi_cross_bar_io_m_port_1_wvalid),
    .io_m_port_1_wready(axi_cross_bar_io_m_port_1_wready),
    .io_m_port_1_bvalid(axi_cross_bar_io_m_port_1_bvalid),
    .io_s_port_arid(axi_cross_bar_io_s_port_arid),
    .io_s_port_araddr(axi_cross_bar_io_s_port_araddr),
    .io_s_port_arlen(axi_cross_bar_io_s_port_arlen),
    .io_s_port_arsize(axi_cross_bar_io_s_port_arsize),
    .io_s_port_arburst(axi_cross_bar_io_s_port_arburst),
    .io_s_port_arvalid(axi_cross_bar_io_s_port_arvalid),
    .io_s_port_arready(axi_cross_bar_io_s_port_arready),
    .io_s_port_rdata(axi_cross_bar_io_s_port_rdata),
    .io_s_port_rlast(axi_cross_bar_io_s_port_rlast),
    .io_s_port_rvalid(axi_cross_bar_io_s_port_rvalid),
    .io_s_port_rready(axi_cross_bar_io_s_port_rready),
    .io_s_port_awid(axi_cross_bar_io_s_port_awid),
    .io_s_port_awaddr(axi_cross_bar_io_s_port_awaddr),
    .io_s_port_awlen(axi_cross_bar_io_s_port_awlen),
    .io_s_port_awsize(axi_cross_bar_io_s_port_awsize),
    .io_s_port_awburst(axi_cross_bar_io_s_port_awburst),
    .io_s_port_awvalid(axi_cross_bar_io_s_port_awvalid),
    .io_s_port_awready(axi_cross_bar_io_s_port_awready),
    .io_s_port_wid(axi_cross_bar_io_s_port_wid),
    .io_s_port_wdata(axi_cross_bar_io_s_port_wdata),
    .io_s_port_wstrb(axi_cross_bar_io_s_port_wstrb),
    .io_s_port_wlast(axi_cross_bar_io_s_port_wlast),
    .io_s_port_wvalid(axi_cross_bar_io_s_port_wvalid),
    .io_s_port_wready(axi_cross_bar_io_s_port_wready),
    .io_s_port_bvalid(axi_cross_bar_io_s_port_bvalid)
  );
  assign io_m_port_0_arready = axi_cross_bar_io_m_port_0_arready; // @[axi_ram_port.scala 205:34]
  assign io_m_port_0_rdata = axi_cross_bar_io_m_port_0_rdata; // @[axi_ram_port.scala 205:34]
  assign io_m_port_0_rlast = axi_cross_bar_io_m_port_0_rlast; // @[axi_ram_port.scala 205:34]
  assign io_m_port_0_rvalid = axi_cross_bar_io_m_port_0_rvalid; // @[axi_ram_port.scala 205:34]
  assign io_m_port_1_arready = axi_cross_bar_io_m_port_1_arready; // @[axi_ram_port.scala 205:34]
  assign io_m_port_1_rdata = axi_cross_bar_io_m_port_1_rdata; // @[axi_ram_port.scala 205:34]
  assign io_m_port_1_rlast = axi_cross_bar_io_m_port_1_rlast; // @[axi_ram_port.scala 205:34]
  assign io_m_port_1_rvalid = axi_cross_bar_io_m_port_1_rvalid; // @[axi_ram_port.scala 205:34]
  assign io_m_port_1_awready = axi_cross_bar_io_m_port_1_awready; // @[axi_ram_port.scala 205:34]
  assign io_m_port_1_wready = axi_cross_bar_io_m_port_1_wready; // @[axi_ram_port.scala 205:34]
  assign io_m_port_1_bvalid = axi_cross_bar_io_m_port_1_bvalid; // @[axi_ram_port.scala 205:34]
  assign io_s_port_0_arid = access_select_s_port_num_r_0 ? axi_cross_bar_io_s_port_arid : 4'h0; // @[axi_ram_port.scala 282:57 283:51 298:51]
  assign io_s_port_0_araddr = access_select_s_port_num_r_0 ? axi_cross_bar_io_s_port_araddr : 64'h0; // @[axi_ram_port.scala 282:57 284:51 299:51]
  assign io_s_port_0_arlen = access_select_s_port_num_r_0 ? axi_cross_bar_io_s_port_arlen : 4'h0; // @[axi_ram_port.scala 282:57 285:51 300:51]
  assign io_s_port_0_arsize = access_select_s_port_num_r_0 ? axi_cross_bar_io_s_port_arsize : 3'h0; // @[axi_ram_port.scala 282:57 286:51 301:51]
  assign io_s_port_0_arburst = access_select_s_port_num_r_0 ? axi_cross_bar_io_s_port_arburst : 2'h0; // @[axi_ram_port.scala 282:57 287:51 302:51]
  assign io_s_port_0_arvalid = access_select_s_port_num_r_0 & axi_cross_bar_io_s_port_arvalid; // @[axi_ram_port.scala 282:57 291:51 306:51]
  assign io_s_port_0_rready = access_select_s_port_num_r_0 & axi_cross_bar_io_s_port_rready; // @[axi_ram_port.scala 282:57 292:51 307:51]
  assign io_s_port_0_awid = access_select_s_port_num_w_0 ? axi_cross_bar_io_s_port_awid : 4'h0; // @[axi_ram_port.scala 309:57 310:52 328:52]
  assign io_s_port_0_awaddr = access_select_s_port_num_w_0 ? axi_cross_bar_io_s_port_awaddr : 64'h0; // @[axi_ram_port.scala 309:57 311:52 329:52]
  assign io_s_port_0_awlen = access_select_s_port_num_w_0 ? axi_cross_bar_io_s_port_awlen : 4'h0; // @[axi_ram_port.scala 309:57 312:52 330:52]
  assign io_s_port_0_awsize = access_select_s_port_num_w_0 ? axi_cross_bar_io_s_port_awsize : 3'h0; // @[axi_ram_port.scala 309:57 313:52 331:52]
  assign io_s_port_0_awburst = access_select_s_port_num_w_0 ? axi_cross_bar_io_s_port_awburst : 2'h0; // @[axi_ram_port.scala 309:57 314:52 332:52]
  assign io_s_port_0_awvalid = access_select_s_port_num_w_0 & axi_cross_bar_io_s_port_awvalid; // @[axi_ram_port.scala 309:57 318:52 336:52]
  assign io_s_port_0_wid = access_select_s_port_num_w_0 ? axi_cross_bar_io_s_port_wid : 4'h0; // @[axi_ram_port.scala 309:57 319:52 337:52]
  assign io_s_port_0_wdata = access_select_s_port_num_w_0 ? axi_cross_bar_io_s_port_wdata : 64'h0; // @[axi_ram_port.scala 309:57 320:52 338:52]
  assign io_s_port_0_wstrb = access_select_s_port_num_w_0 ? axi_cross_bar_io_s_port_wstrb : 8'h0; // @[axi_ram_port.scala 309:57 321:52 339:52]
  assign io_s_port_0_wlast = access_select_s_port_num_w_0 & axi_cross_bar_io_s_port_wlast; // @[axi_ram_port.scala 309:57 322:52 340:52]
  assign io_s_port_0_wvalid = access_select_s_port_num_w_0 & axi_cross_bar_io_s_port_wvalid; // @[axi_ram_port.scala 309:57 323:52 341:52]
  assign io_s_port_0_bready = access_select_s_port_num_w_0 & axi_cross_bar_io_s_port_bvalid; // @[axi_ram_port.scala 309:57 324:52 342:52]
  assign io_s_port_1_araddr = access_select_s_port_num_r_1 ? axi_cross_bar_io_s_port_araddr : 64'h0; // @[axi_ram_port.scala 282:57 284:51 299:51]
  assign io_s_port_1_arvalid = access_select_s_port_num_r_1 & axi_cross_bar_io_s_port_arvalid; // @[axi_ram_port.scala 282:57 291:51 306:51]
  assign io_s_port_1_rready = access_select_s_port_num_r_1 & axi_cross_bar_io_s_port_rready; // @[axi_ram_port.scala 282:57 292:51 307:51]
  assign io_s_port_1_awaddr = access_select_s_port_num_w_1 ? axi_cross_bar_io_s_port_awaddr : 64'h0; // @[axi_ram_port.scala 309:57 311:52 329:52]
  assign io_s_port_1_awsize = access_select_s_port_num_w_1 ? axi_cross_bar_io_s_port_awsize : 3'h0; // @[axi_ram_port.scala 309:57 313:52 331:52]
  assign io_s_port_1_awvalid = access_select_s_port_num_w_1 & axi_cross_bar_io_s_port_awvalid; // @[axi_ram_port.scala 309:57 318:52 336:52]
  assign io_s_port_1_wdata = access_select_s_port_num_w_1 ? axi_cross_bar_io_s_port_wdata : 64'h0; // @[axi_ram_port.scala 309:57 320:52 338:52]
  assign io_s_port_1_wvalid = access_select_s_port_num_w_1 & axi_cross_bar_io_s_port_wvalid; // @[axi_ram_port.scala 309:57 323:52 341:52]
  assign axi_cross_bar_clock = clock;
  assign axi_cross_bar_reset = reset;
  assign axi_cross_bar_io_m_port_0_araddr = io_m_port_0_araddr; // @[axi_ram_port.scala 205:34]
  assign axi_cross_bar_io_m_port_0_arlen = io_m_port_0_arlen; // @[axi_ram_port.scala 205:34]
  assign axi_cross_bar_io_m_port_0_arburst = io_m_port_0_arburst; // @[axi_ram_port.scala 205:34]
  assign axi_cross_bar_io_m_port_0_arvalid = io_m_port_0_arvalid; // @[axi_ram_port.scala 205:34]
  assign axi_cross_bar_io_m_port_1_araddr = io_m_port_1_araddr; // @[axi_ram_port.scala 205:34]
  assign axi_cross_bar_io_m_port_1_arlen = io_m_port_1_arlen; // @[axi_ram_port.scala 205:34]
  assign axi_cross_bar_io_m_port_1_arsize = io_m_port_1_arsize; // @[axi_ram_port.scala 205:34]
  assign axi_cross_bar_io_m_port_1_arburst = io_m_port_1_arburst; // @[axi_ram_port.scala 205:34]
  assign axi_cross_bar_io_m_port_1_arvalid = io_m_port_1_arvalid; // @[axi_ram_port.scala 205:34]
  assign axi_cross_bar_io_m_port_1_awaddr = io_m_port_1_awaddr; // @[axi_ram_port.scala 205:34]
  assign axi_cross_bar_io_m_port_1_awlen = io_m_port_1_awlen; // @[axi_ram_port.scala 205:34]
  assign axi_cross_bar_io_m_port_1_awsize = io_m_port_1_awsize; // @[axi_ram_port.scala 205:34]
  assign axi_cross_bar_io_m_port_1_awburst = io_m_port_1_awburst; // @[axi_ram_port.scala 205:34]
  assign axi_cross_bar_io_m_port_1_awvalid = io_m_port_1_awvalid; // @[axi_ram_port.scala 205:34]
  assign axi_cross_bar_io_m_port_1_wdata = io_m_port_1_wdata; // @[axi_ram_port.scala 205:34]
  assign axi_cross_bar_io_m_port_1_wstrb = io_m_port_1_wstrb; // @[axi_ram_port.scala 205:34]
  assign axi_cross_bar_io_m_port_1_wlast = io_m_port_1_wlast; // @[axi_ram_port.scala 205:34]
  assign axi_cross_bar_io_m_port_1_wvalid = io_m_port_1_wvalid; // @[axi_ram_port.scala 205:34]
  assign axi_cross_bar_io_s_port_arready = _T_17[0]; // @[axi_ram_port.scala 353:49]
  assign axi_cross_bar_io_s_port_rdata = _T_21 | _T_22; // @[Mux.scala 27:73]
  assign axi_cross_bar_io_s_port_rlast = access_select_s_port_num_r_0 & io_s_port_0_rlast | access_select_s_port_num_r_1
     & io_s_port_1_rlast; // @[Mux.scala 27:73]
  assign axi_cross_bar_io_s_port_rvalid = access_select_s_port_num_r_0 & io_s_port_0_rvalid |
    access_select_s_port_num_r_1 & io_s_port_1_rvalid; // @[Mux.scala 27:73]
  assign axi_cross_bar_io_s_port_awready = access_select_s_port_num_w_0 & io_s_port_0_awready |
    access_select_s_port_num_w_1; // @[Mux.scala 27:73]
  assign axi_cross_bar_io_s_port_wready = access_select_s_port_num_w_0 & io_s_port_0_wready |
    access_select_s_port_num_w_1 & io_s_port_1_wready; // @[Mux.scala 27:73]
  assign axi_cross_bar_io_s_port_bvalid = access_select_s_port_num_w_0 & io_s_port_0_bvalid |
    access_select_s_port_num_w_1 & io_s_port_1_bvalid; // @[Mux.scala 27:73]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[axi_ram_port.scala 217:50]
      select_s_port_num_r_0 <= 1'h0;
    end else if (_r_to_be_T[1]) begin
      select_s_port_num_r_0 <= 1'h0;
    end else begin
      select_s_port_num_r_0 <= 1'h1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[axi_ram_port.scala 234:42]
      select_s_port_num_r_1 <= 1'h0;
    end else if (_access_select_s_port_num_r_1_T) begin // @[axi_ram_port.scala 235:108]
      select_s_port_num_r_1 <= _access_select_s_port_num_r_1_T_3;
    end else if (io_s_port_1_rlast) begin
      select_s_port_num_r_1 <= 1'h0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[axi_ram_port.scala 221:50]
      select_s_port_num_w_0 <= 1'h0;
    end else if (_w_to_be_T[1]) begin
      select_s_port_num_w_0 <= 1'h0;
    end else begin
      select_s_port_num_w_0 <= 1'h1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[axi_ram_port.scala 239:42]
      select_s_port_num_w_1 <= 1'h0;
    end else if (_access_select_s_port_num_w_1_T) begin // @[axi_ram_port.scala 240:108]
      select_s_port_num_w_1 <= _access_select_s_port_num_w_1_T_3;
    end else if (io_s_port_1_bvalid) begin
      select_s_port_num_w_1 <= 1'h0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  select_s_port_num_r_0 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  select_s_port_num_r_1 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  select_s_port_num_w_0 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  select_s_port_num_w_1 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    select_s_port_num_r_0 = 1'h0;
  end
  if (reset) begin
    select_s_port_num_r_1 = 1'h0;
  end
  if (reset) begin
    select_s_port_num_w_0 = 1'h0;
  end
  if (reset) begin
    select_s_port_num_w_1 = 1'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module timer_periph(
  input         clock,
  input         reset,
  input  [63:0] io_axi_port_araddr,
  input         io_axi_port_arvalid,
  output        io_axi_port_arready,
  output [63:0] io_axi_port_rdata,
  output        io_axi_port_rlast,
  output        io_axi_port_rvalid,
  input         io_axi_port_rready,
  input  [63:0] io_axi_port_awaddr,
  input  [2:0]  io_axi_port_awsize,
  input         io_axi_port_awvalid,
  output        io_axi_port_awready,
  input  [63:0] io_axi_port_wdata,
  input         io_axi_port_wvalid,
  output        io_axi_port_wready,
  output        io_axi_port_bvalid,
  output        io_int_line
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtime; // @[clint.scala 25:26]
  reg [63:0] mtimecmp; // @[clint.scala 26:27]
  reg [31:0] msip; // @[clint.scala 27:25]
  reg [2:0] axi_read_state; // @[clint.scala 30:33]
  reg [2:0] axi_write_state; // @[clint.scala 31:34]
  reg [63:0] axi_read_addr; // @[clint.scala 32:32]
  reg [63:0] axi_write_addr; // @[clint.scala 33:33]
  reg [3:0] axi_write_size; // @[clint.scala 34:33]
  wire  _axi_read_state_T_2 = io_axi_port_arvalid & io_axi_port_arready; // @[clint.scala 38:54]
  wire  _axi_write_state_T_2 = io_axi_port_awvalid & io_axi_port_awready; // @[clint.scala 43:54]
  wire [1:0] _axi_write_size_T_6 = 3'h1 == io_axi_port_awsize ? 2'h2 : {{1'd0}, 3'h0 == io_axi_port_awsize}; // @[Mux.scala 81:58]
  wire [2:0] _axi_write_size_T_8 = 3'h2 == io_axi_port_awsize ? 3'h4 : {{1'd0}, _axi_write_size_T_6}; // @[Mux.scala 81:58]
  wire [5:0] _axi_write_data_T_1 = {io_axi_port_awaddr[2:0], 3'h0}; // @[clint.scala 51:69]
  wire [126:0] _GEN_0 = {{63'd0}, io_axi_port_wdata}; // @[clint.scala 51:41]
  wire [126:0] _axi_write_data_T_2 = _GEN_0 << _axi_write_data_T_1; // @[clint.scala 51:41]
  wire [31:0] _read_data_T_7 = 64'h20000000 == axi_read_addr ? msip : 32'h0; // @[Mux.scala 81:58]
  wire [63:0] _read_data_T_9 = 64'h2000bff8 == axi_read_addr ? mtime : {{32'd0}, _read_data_T_7}; // @[Mux.scala 81:58]
  wire [3:0] _mtime_to_be_0_T_3 = {1'h0,axi_write_addr[2:0]}; // @[Cat.scala 31:58]
  wire [3:0] _mtime_to_be_0_T_5 = _mtime_to_be_0_T_3 + axi_write_size; // @[clint.scala 70:109]
  wire  _mtime_to_be_0_T_7 = axi_write_addr[2:0] <= 3'h0 & _mtime_to_be_0_T_5 > 4'h0; // @[clint.scala 70:70]
  wire [63:0] axi_write_data = _axi_write_data_T_2[63:0]; // @[clint.scala 35:30 51:20]
  wire [7:0] mtime_to_be_0 = axi_write_addr[2:0] <= 3'h0 & _mtime_to_be_0_T_5 > 4'h0 ? axi_write_data[7:0] : mtime[7:0]; // @[clint.scala 70:38]
  wire  _mtime_to_be_1_T_7 = axi_write_addr[2:0] <= 3'h1 & _mtime_to_be_0_T_5 > 4'h1; // @[clint.scala 70:70]
  wire [7:0] mtime_to_be_1 = axi_write_addr[2:0] <= 3'h1 & _mtime_to_be_0_T_5 > 4'h1 ? axi_write_data[15:8] : mtime[15:8
    ]; // @[clint.scala 70:38]
  wire  _mtime_to_be_2_T_7 = axi_write_addr[2:0] <= 3'h2 & _mtime_to_be_0_T_5 > 4'h2; // @[clint.scala 70:70]
  wire [7:0] mtime_to_be_2 = axi_write_addr[2:0] <= 3'h2 & _mtime_to_be_0_T_5 > 4'h2 ? axi_write_data[23:16] : mtime[23:
    16]; // @[clint.scala 70:38]
  wire  _mtime_to_be_3_T_7 = axi_write_addr[2:0] <= 3'h3 & _mtime_to_be_0_T_5 > 4'h3; // @[clint.scala 70:70]
  wire [7:0] mtime_to_be_3 = axi_write_addr[2:0] <= 3'h3 & _mtime_to_be_0_T_5 > 4'h3 ? axi_write_data[31:24] : mtime[31:
    24]; // @[clint.scala 70:38]
  wire  _mtime_to_be_4_T_7 = axi_write_addr[2:0] <= 3'h4 & _mtime_to_be_0_T_5 > 4'h4; // @[clint.scala 70:70]
  wire [7:0] mtime_to_be_4 = axi_write_addr[2:0] <= 3'h4 & _mtime_to_be_0_T_5 > 4'h4 ? axi_write_data[39:32] : mtime[39:
    32]; // @[clint.scala 70:38]
  wire  _mtime_to_be_5_T_7 = axi_write_addr[2:0] <= 3'h5 & _mtime_to_be_0_T_5 > 4'h5; // @[clint.scala 70:70]
  wire [7:0] mtime_to_be_5 = axi_write_addr[2:0] <= 3'h5 & _mtime_to_be_0_T_5 > 4'h5 ? axi_write_data[47:40] : mtime[47:
    40]; // @[clint.scala 70:38]
  wire  _mtime_to_be_6_T_7 = axi_write_addr[2:0] <= 3'h6 & _mtime_to_be_0_T_5 > 4'h6; // @[clint.scala 70:70]
  wire [7:0] mtime_to_be_6 = axi_write_addr[2:0] <= 3'h6 & _mtime_to_be_0_T_5 > 4'h6 ? axi_write_data[55:48] : mtime[55:
    48]; // @[clint.scala 70:38]
  wire  _mtime_to_be_7_T_6 = _mtime_to_be_0_T_5 > 4'h7; // @[clint.scala 70:126]
  wire [7:0] mtime_to_be_7 = _mtime_to_be_0_T_5 > 4'h7 ? axi_write_data[63:56] : mtime[63:56]; // @[clint.scala 70:38]
  wire  _mtime_T_2 = axi_write_state == 3'h1 & io_axi_port_wvalid; // @[clint.scala 73:48]
  wire [63:0] _mtime_T_9 = {mtime_to_be_7,mtime_to_be_6,mtime_to_be_5,mtime_to_be_4,mtime_to_be_3,mtime_to_be_2,
    mtime_to_be_1,mtime_to_be_0}; // @[clint.scala 74:21]
  wire [63:0] _mtime_T_11 = mtime + 64'h1; // @[clint.scala 74:34]
  wire [7:0] mtimecmp_to_be_0 = _mtime_to_be_0_T_7 ? axi_write_data[7:0] : mtimecmp[7:0]; // @[clint.scala 77:41]
  wire [7:0] mtimecmp_to_be_1 = _mtime_to_be_1_T_7 ? axi_write_data[15:8] : mtimecmp[15:8]; // @[clint.scala 77:41]
  wire [7:0] mtimecmp_to_be_2 = _mtime_to_be_2_T_7 ? axi_write_data[23:16] : mtimecmp[23:16]; // @[clint.scala 77:41]
  wire [7:0] mtimecmp_to_be_3 = _mtime_to_be_3_T_7 ? axi_write_data[31:24] : mtimecmp[31:24]; // @[clint.scala 77:41]
  wire [7:0] mtimecmp_to_be_4 = _mtime_to_be_4_T_7 ? axi_write_data[39:32] : mtimecmp[39:32]; // @[clint.scala 77:41]
  wire [7:0] mtimecmp_to_be_5 = _mtime_to_be_5_T_7 ? axi_write_data[47:40] : mtimecmp[47:40]; // @[clint.scala 77:41]
  wire [7:0] mtimecmp_to_be_6 = _mtime_to_be_6_T_7 ? axi_write_data[55:48] : mtimecmp[55:48]; // @[clint.scala 77:41]
  wire [7:0] mtimecmp_to_be_7 = _mtime_to_be_7_T_6 ? axi_write_data[63:56] : mtimecmp[63:56]; // @[clint.scala 77:41]
  wire [63:0] _mtimecmp_T_9 = {mtimecmp_to_be_7,mtimecmp_to_be_6,mtimecmp_to_be_5,mtimecmp_to_be_4,mtimecmp_to_be_3,
    mtimecmp_to_be_2,mtimecmp_to_be_1,mtimecmp_to_be_0}; // @[clint.scala 81:24]
  wire [31:0] _msip_T_8 = {31'h0,axi_write_data[0]}; // @[Cat.scala 31:58]
  assign io_axi_port_arready = 1'h1; // @[clint.scala 63:25]
  assign io_axi_port_rdata = 64'h20004000 == axi_read_addr ? mtimecmp : _read_data_T_9; // @[Mux.scala 81:58]
  assign io_axi_port_rlast = axi_read_state == 3'h1 & io_axi_port_rready; // @[clint.scala 61:55]
  assign io_axi_port_rvalid = axi_read_state == 3'h1; // @[clint.scala 62:42]
  assign io_axi_port_awready = 1'h1; // @[clint.scala 85:26]
  assign io_axi_port_wready = axi_write_state == 3'h1; // @[clint.scala 86:45]
  assign io_axi_port_bvalid = axi_write_state == 3'h2; // @[clint.scala 89:45]
  assign io_int_line = mtime >= mtimecmp; // @[clint.scala 91:26]
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[clint.scala 73:17]
      mtime <= 64'h0;
    end else if (axi_write_state == 3'h1 & io_axi_port_wvalid & axi_write_addr[63:3] == 61'h40017ff) begin
      mtime <= _mtime_T_9;
    end else begin
      mtime <= _mtime_T_11;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[clint.scala 80:20]
      mtimecmp <= 64'h0;
    end else if (_mtime_T_2 & axi_write_addr[63:3] == 61'h4000800) begin
      mtimecmp <= _mtimecmp_T_9;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[clint.scala 82:16]
      msip <= 32'h0;
    end else if (axi_read_addr == 64'h1 & io_axi_port_wvalid & axi_write_addr == 64'h20000000) begin
      msip <= _msip_T_8;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Mux.scala 81:58]
      axi_read_state <= 3'h0; // @[clint.scala 39:26]
    end else if (3'h1 == axi_read_state) begin // @[Mux.scala 81:58]
      if (!(io_axi_port_rready)) begin // @[clint.scala 38:26]
        axi_read_state <= 3'h0;
      end
    end else if (3'h0 == axi_read_state) begin
      if (io_axi_port_arvalid & io_axi_port_arready) begin
        axi_read_state <= 3'h1;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[Mux.scala 81:58]
      axi_write_state <= 3'h0;
    end else if (3'h2 == axi_write_state) begin // @[Mux.scala 81:58]
      axi_write_state <= 3'h0; // @[clint.scala 44:26]
    end else if (3'h1 == axi_write_state) begin // @[Mux.scala 81:58]
      if (io_axi_port_wready) begin // @[clint.scala 43:26]
        axi_write_state <= 3'h2;
      end
    end else if (3'h0 == axi_write_state) begin
      if (io_axi_port_awvalid & io_axi_port_awready) begin
        axi_write_state <= 3'h1;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[clint.scala 48:25]
      axi_read_addr <= 64'h0;
    end else if (_axi_read_state_T_2) begin
      axi_read_addr <= io_axi_port_araddr;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[clint.scala 49:26]
      axi_write_addr <= 64'h0;
    end else if (_axi_write_state_T_2) begin
      axi_write_addr <= io_axi_port_awaddr;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin // @[clint.scala 50:26]
      axi_write_size <= 4'h0; // @[Mux.scala 81:58]
    end else if (_axi_write_state_T_2) begin
      if (3'h3 == io_axi_port_awsize) begin
        axi_write_size <= 4'h8;
      end else begin
        axi_write_size <= {{1'd0}, _axi_write_size_T_8};
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtime = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mtimecmp = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  msip = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  axi_read_state = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  axi_write_state = _RAND_4[2:0];
  _RAND_5 = {2{`RANDOM}};
  axi_read_addr = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  axi_write_addr = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  axi_write_size = _RAND_7[3:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    mtime = 64'h0;
  end
  if (reset) begin
    mtimecmp = 64'h0;
  end
  if (reset) begin
    msip = 32'h0;
  end
  if (reset) begin
    axi_read_state = 3'h0;
  end
  if (reset) begin
    axi_write_state = 3'h0;
  end
  if (reset) begin
    axi_read_addr = 64'h0;
  end
  if (reset) begin
    axi_write_addr = 64'h0;
  end
  if (reset) begin
    axi_write_size = 4'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module mycpu_top(
  input         aresetn,
  input         aclk,
  output [3:0]  axi_mem_port_arid,
  output [63:0] axi_mem_port_araddr,
  output [3:0]  axi_mem_port_arlen,
  output [2:0]  axi_mem_port_arsize,
  output [1:0]  axi_mem_port_arburst,
  output [1:0]  axi_mem_port_arlock,
  output [3:0]  axi_mem_port_arcache,
  output [2:0]  axi_mem_port_arprot,
  output        axi_mem_port_arvalid,
  input         axi_mem_port_arready,
  input  [3:0]  axi_mem_port_rid,
  input  [63:0] axi_mem_port_rdata,
  input  [1:0]  axi_mem_port_rresp,
  input         axi_mem_port_rlast,
  input         axi_mem_port_rvalid,
  output        axi_mem_port_rready,
  output [3:0]  axi_mem_port_awid,
  output [63:0] axi_mem_port_awaddr,
  output [3:0]  axi_mem_port_awlen,
  output [2:0]  axi_mem_port_awsize,
  output [1:0]  axi_mem_port_awburst,
  output [1:0]  axi_mem_port_awlock,
  output [3:0]  axi_mem_port_awcache,
  output [2:0]  axi_mem_port_awprot,
  output        axi_mem_port_awvalid,
  input         axi_mem_port_awready,
  output [3:0]  axi_mem_port_wid,
  output [63:0] axi_mem_port_wdata,
  output [7:0]  axi_mem_port_wstrb,
  output        axi_mem_port_wlast,
  output        axi_mem_port_wvalid,
  input         axi_mem_port_wready,
  input  [3:0]  axi_mem_port_bid,
  input  [1:0]  axi_mem_port_bresp,
  input         axi_mem_port_bvalid,
  output        axi_mem_port_bready,
  output [31:0] debug_wb_pc,
  output [3:0]  debug_wb_rf_wen,
  output [4:0]  debug_wb_rf_wnum,
  output [31:0] debug_wb_rf_wdata
);
  wire  u_riscv_cpu_ext_int_timer; // @[my_cpu_top.scala 127:29]
  wire  u_riscv_cpu_resetn; // @[my_cpu_top.scala 127:29]
  wire  u_riscv_cpu_clk; // @[my_cpu_top.scala 127:29]
  wire  u_riscv_cpu_inst_cache; // @[my_cpu_top.scala 127:29]
  wire  u_riscv_cpu_inst_sram_en; // @[my_cpu_top.scala 127:29]
  wire [63:0] u_riscv_cpu_inst_sram_addr; // @[my_cpu_top.scala 127:29]
  wire [39:0] u_riscv_cpu_inst_sram_rdata_L; // @[my_cpu_top.scala 127:29]
  wire [1:0] u_riscv_cpu_inst_write_en; // @[my_cpu_top.scala 127:29]
  wire  u_riscv_cpu_stage2_flush; // @[my_cpu_top.scala 127:29]
  wire  u_riscv_cpu_stage2_stall; // @[my_cpu_top.scala 127:29]
  wire  u_riscv_cpu_stage1_valid_flush; // @[my_cpu_top.scala 127:29]
  wire  u_riscv_cpu_inst_ready_to_use; // @[my_cpu_top.scala 127:29]
  wire  u_riscv_cpu_inst_buffer_full; // @[my_cpu_top.scala 127:29]
  wire  u_riscv_cpu_data_sram_en; // @[my_cpu_top.scala 127:29]
  wire  u_riscv_cpu_data_sram_wen; // @[my_cpu_top.scala 127:29]
  wire [1:0] u_riscv_cpu_data_size; // @[my_cpu_top.scala 127:29]
  wire [63:0] u_riscv_cpu_data_sram_addr; // @[my_cpu_top.scala 127:29]
  wire [63:0] u_riscv_cpu_data_sram_wdata; // @[my_cpu_top.scala 127:29]
  wire  u_riscv_cpu_data_cache; // @[my_cpu_top.scala 127:29]
  wire [63:0] u_riscv_cpu_data_sram_rdata; // @[my_cpu_top.scala 127:29]
  wire  u_riscv_cpu_data_stage2_stall; // @[my_cpu_top.scala 127:29]
  wire [7:0] u_riscv_cpu_data_wstrb; // @[my_cpu_top.scala 127:29]
  wire  u_riscv_cpu_data_fence_i_control; // @[my_cpu_top.scala 127:29]
  wire [63:0] u_riscv_cpu_debug_wb_pc; // @[my_cpu_top.scala 127:29]
  wire [3:0] u_riscv_cpu_debug_wb_rf_wen; // @[my_cpu_top.scala 127:29]
  wire [4:0] u_riscv_cpu_debug_wb_rf_wnum; // @[my_cpu_top.scala 127:29]
  wire [63:0] u_riscv_cpu_debug_wb_rf_wdata; // @[my_cpu_top.scala 127:29]
  wire  u_riscv_cpu_icache_tag_flush; // @[my_cpu_top.scala 127:29]
  wire  inst_cache_clock; // @[my_cpu_top.scala 128:30]
  wire  inst_cache_reset; // @[my_cpu_top.scala 128:30]
  wire [63:0] inst_cache_io_port_araddr; // @[my_cpu_top.scala 128:30]
  wire [3:0] inst_cache_io_port_arlen; // @[my_cpu_top.scala 128:30]
  wire [1:0] inst_cache_io_port_arburst; // @[my_cpu_top.scala 128:30]
  wire  inst_cache_io_port_arvalid; // @[my_cpu_top.scala 128:30]
  wire  inst_cache_io_port_arready; // @[my_cpu_top.scala 128:30]
  wire [63:0] inst_cache_io_port_rdata; // @[my_cpu_top.scala 128:30]
  wire  inst_cache_io_port_rlast; // @[my_cpu_top.scala 128:30]
  wire  inst_cache_io_port_rvalid; // @[my_cpu_top.scala 128:30]
  wire  inst_cache_io_stage2_flush; // @[my_cpu_top.scala 128:30]
  wire  inst_cache_io_stage2_stall; // @[my_cpu_top.scala 128:30]
  wire  inst_cache_io_stage1_valid_flush; // @[my_cpu_top.scala 128:30]
  wire  inst_cache_io_inst_ready_to_use; // @[my_cpu_top.scala 128:30]
  wire  inst_cache_io_inst_buffer_full; // @[my_cpu_top.scala 128:30]
  wire [63:0] inst_cache_io_v_addr_for_tlb; // @[my_cpu_top.scala 128:30]
  wire [63:0] inst_cache_io_p_addr_for_tlb; // @[my_cpu_top.scala 128:30]
  wire  inst_cache_io_sram_req; // @[my_cpu_top.scala 128:30]
  wire [63:0] inst_cache_io_sram_addr; // @[my_cpu_top.scala 128:30]
  wire [1:0] inst_cache_io_sram_write_en; // @[my_cpu_top.scala 128:30]
  wire [39:0] inst_cache_io_sram_rdata_L; // @[my_cpu_top.scala 128:30]
  wire  inst_cache_io_sram_cache; // @[my_cpu_top.scala 128:30]
  wire  inst_cache_io_tag_valid_flush; // @[my_cpu_top.scala 128:30]
  wire  data_cache_clock; // @[my_cpu_top.scala 130:30]
  wire  data_cache_reset; // @[my_cpu_top.scala 130:30]
  wire [63:0] data_cache_io_port_araddr; // @[my_cpu_top.scala 130:30]
  wire [3:0] data_cache_io_port_arlen; // @[my_cpu_top.scala 130:30]
  wire [2:0] data_cache_io_port_arsize; // @[my_cpu_top.scala 130:30]
  wire [1:0] data_cache_io_port_arburst; // @[my_cpu_top.scala 130:30]
  wire  data_cache_io_port_arvalid; // @[my_cpu_top.scala 130:30]
  wire  data_cache_io_port_arready; // @[my_cpu_top.scala 130:30]
  wire [63:0] data_cache_io_port_rdata; // @[my_cpu_top.scala 130:30]
  wire  data_cache_io_port_rlast; // @[my_cpu_top.scala 130:30]
  wire  data_cache_io_port_rvalid; // @[my_cpu_top.scala 130:30]
  wire [63:0] data_cache_io_port_awaddr; // @[my_cpu_top.scala 130:30]
  wire [3:0] data_cache_io_port_awlen; // @[my_cpu_top.scala 130:30]
  wire [2:0] data_cache_io_port_awsize; // @[my_cpu_top.scala 130:30]
  wire [1:0] data_cache_io_port_awburst; // @[my_cpu_top.scala 130:30]
  wire  data_cache_io_port_awvalid; // @[my_cpu_top.scala 130:30]
  wire  data_cache_io_port_awready; // @[my_cpu_top.scala 130:30]
  wire [63:0] data_cache_io_port_wdata; // @[my_cpu_top.scala 130:30]
  wire [7:0] data_cache_io_port_wstrb; // @[my_cpu_top.scala 130:30]
  wire  data_cache_io_port_wlast; // @[my_cpu_top.scala 130:30]
  wire  data_cache_io_port_wvalid; // @[my_cpu_top.scala 130:30]
  wire  data_cache_io_port_wready; // @[my_cpu_top.scala 130:30]
  wire  data_cache_io_port_bvalid; // @[my_cpu_top.scala 130:30]
  wire  data_cache_io_stage2_stall; // @[my_cpu_top.scala 130:30]
  wire [63:0] data_cache_io_v_addr_for_tlb; // @[my_cpu_top.scala 130:30]
  wire [63:0] data_cache_io_p_addr_for_tlb; // @[my_cpu_top.scala 130:30]
  wire  data_cache_io_tlb_req; // @[my_cpu_top.scala 130:30]
  wire [7:0] data_cache_io_data_wstrb; // @[my_cpu_top.scala 130:30]
  wire  data_cache_io_sram_req; // @[my_cpu_top.scala 130:30]
  wire  data_cache_io_sram_wr; // @[my_cpu_top.scala 130:30]
  wire [2:0] data_cache_io_sram_size; // @[my_cpu_top.scala 130:30]
  wire [63:0] data_cache_io_sram_addr; // @[my_cpu_top.scala 130:30]
  wire [63:0] data_cache_io_sram_wdata; // @[my_cpu_top.scala 130:30]
  wire [63:0] data_cache_io_sram_rdata; // @[my_cpu_top.scala 130:30]
  wire  data_cache_io_sram_cache; // @[my_cpu_top.scala 130:30]
  wire  data_cache_io_fence_i_control; // @[my_cpu_top.scala 130:30]
  wire  _axi_cross_bar_clock; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_reset; // @[my_cpu_top.scala 132:32]
  wire [63:0] _axi_cross_bar_io_m_port_0_araddr; // @[my_cpu_top.scala 132:32]
  wire [3:0] _axi_cross_bar_io_m_port_0_arlen; // @[my_cpu_top.scala 132:32]
  wire [1:0] _axi_cross_bar_io_m_port_0_arburst; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_m_port_0_arvalid; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_m_port_0_arready; // @[my_cpu_top.scala 132:32]
  wire [63:0] _axi_cross_bar_io_m_port_0_rdata; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_m_port_0_rlast; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_m_port_0_rvalid; // @[my_cpu_top.scala 132:32]
  wire [63:0] _axi_cross_bar_io_m_port_1_araddr; // @[my_cpu_top.scala 132:32]
  wire [3:0] _axi_cross_bar_io_m_port_1_arlen; // @[my_cpu_top.scala 132:32]
  wire [2:0] _axi_cross_bar_io_m_port_1_arsize; // @[my_cpu_top.scala 132:32]
  wire [1:0] _axi_cross_bar_io_m_port_1_arburst; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_m_port_1_arvalid; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_m_port_1_arready; // @[my_cpu_top.scala 132:32]
  wire [63:0] _axi_cross_bar_io_m_port_1_rdata; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_m_port_1_rlast; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_m_port_1_rvalid; // @[my_cpu_top.scala 132:32]
  wire [63:0] _axi_cross_bar_io_m_port_1_awaddr; // @[my_cpu_top.scala 132:32]
  wire [3:0] _axi_cross_bar_io_m_port_1_awlen; // @[my_cpu_top.scala 132:32]
  wire [2:0] _axi_cross_bar_io_m_port_1_awsize; // @[my_cpu_top.scala 132:32]
  wire [1:0] _axi_cross_bar_io_m_port_1_awburst; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_m_port_1_awvalid; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_m_port_1_awready; // @[my_cpu_top.scala 132:32]
  wire [63:0] _axi_cross_bar_io_m_port_1_wdata; // @[my_cpu_top.scala 132:32]
  wire [7:0] _axi_cross_bar_io_m_port_1_wstrb; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_m_port_1_wlast; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_m_port_1_wvalid; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_m_port_1_wready; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_m_port_1_bvalid; // @[my_cpu_top.scala 132:32]
  wire [3:0] _axi_cross_bar_io_s_port_0_arid; // @[my_cpu_top.scala 132:32]
  wire [63:0] _axi_cross_bar_io_s_port_0_araddr; // @[my_cpu_top.scala 132:32]
  wire [3:0] _axi_cross_bar_io_s_port_0_arlen; // @[my_cpu_top.scala 132:32]
  wire [2:0] _axi_cross_bar_io_s_port_0_arsize; // @[my_cpu_top.scala 132:32]
  wire [1:0] _axi_cross_bar_io_s_port_0_arburst; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_s_port_0_arvalid; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_s_port_0_arready; // @[my_cpu_top.scala 132:32]
  wire [63:0] _axi_cross_bar_io_s_port_0_rdata; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_s_port_0_rlast; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_s_port_0_rvalid; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_s_port_0_rready; // @[my_cpu_top.scala 132:32]
  wire [3:0] _axi_cross_bar_io_s_port_0_awid; // @[my_cpu_top.scala 132:32]
  wire [63:0] _axi_cross_bar_io_s_port_0_awaddr; // @[my_cpu_top.scala 132:32]
  wire [3:0] _axi_cross_bar_io_s_port_0_awlen; // @[my_cpu_top.scala 132:32]
  wire [2:0] _axi_cross_bar_io_s_port_0_awsize; // @[my_cpu_top.scala 132:32]
  wire [1:0] _axi_cross_bar_io_s_port_0_awburst; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_s_port_0_awvalid; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_s_port_0_awready; // @[my_cpu_top.scala 132:32]
  wire [3:0] _axi_cross_bar_io_s_port_0_wid; // @[my_cpu_top.scala 132:32]
  wire [63:0] _axi_cross_bar_io_s_port_0_wdata; // @[my_cpu_top.scala 132:32]
  wire [7:0] _axi_cross_bar_io_s_port_0_wstrb; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_s_port_0_wlast; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_s_port_0_wvalid; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_s_port_0_wready; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_s_port_0_bvalid; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_s_port_0_bready; // @[my_cpu_top.scala 132:32]
  wire [63:0] _axi_cross_bar_io_s_port_1_araddr; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_s_port_1_arvalid; // @[my_cpu_top.scala 132:32]
  wire [63:0] _axi_cross_bar_io_s_port_1_rdata; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_s_port_1_rlast; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_s_port_1_rvalid; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_s_port_1_rready; // @[my_cpu_top.scala 132:32]
  wire [63:0] _axi_cross_bar_io_s_port_1_awaddr; // @[my_cpu_top.scala 132:32]
  wire [2:0] _axi_cross_bar_io_s_port_1_awsize; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_s_port_1_awvalid; // @[my_cpu_top.scala 132:32]
  wire [63:0] _axi_cross_bar_io_s_port_1_wdata; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_s_port_1_wvalid; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_s_port_1_wready; // @[my_cpu_top.scala 132:32]
  wire  _axi_cross_bar_io_s_port_1_bvalid; // @[my_cpu_top.scala 132:32]
  wire  timer_periph_clock; // @[my_cpu_top.scala 242:27]
  wire  timer_periph_reset; // @[my_cpu_top.scala 242:27]
  wire [63:0] timer_periph_io_axi_port_araddr; // @[my_cpu_top.scala 242:27]
  wire  timer_periph_io_axi_port_arvalid; // @[my_cpu_top.scala 242:27]
  wire  timer_periph_io_axi_port_arready; // @[my_cpu_top.scala 242:27]
  wire [63:0] timer_periph_io_axi_port_rdata; // @[my_cpu_top.scala 242:27]
  wire  timer_periph_io_axi_port_rlast; // @[my_cpu_top.scala 242:27]
  wire  timer_periph_io_axi_port_rvalid; // @[my_cpu_top.scala 242:27]
  wire  timer_periph_io_axi_port_rready; // @[my_cpu_top.scala 242:27]
  wire [63:0] timer_periph_io_axi_port_awaddr; // @[my_cpu_top.scala 242:27]
  wire [2:0] timer_periph_io_axi_port_awsize; // @[my_cpu_top.scala 242:27]
  wire  timer_periph_io_axi_port_awvalid; // @[my_cpu_top.scala 242:27]
  wire  timer_periph_io_axi_port_awready; // @[my_cpu_top.scala 242:27]
  wire [63:0] timer_periph_io_axi_port_wdata; // @[my_cpu_top.scala 242:27]
  wire  timer_periph_io_axi_port_wvalid; // @[my_cpu_top.scala 242:27]
  wire  timer_periph_io_axi_port_wready; // @[my_cpu_top.scala 242:27]
  wire  timer_periph_io_axi_port_bvalid; // @[my_cpu_top.scala 242:27]
  wire  timer_periph_io_int_line; // @[my_cpu_top.scala 242:27]
  myCPU u_riscv_cpu ( // @[my_cpu_top.scala 127:29]
    .ext_int_timer(u_riscv_cpu_ext_int_timer),
    .resetn(u_riscv_cpu_resetn),
    .clk(u_riscv_cpu_clk),
    .inst_cache(u_riscv_cpu_inst_cache),
    .inst_sram_en(u_riscv_cpu_inst_sram_en),
    .inst_sram_addr(u_riscv_cpu_inst_sram_addr),
    .inst_sram_rdata_L(u_riscv_cpu_inst_sram_rdata_L),
    .inst_write_en(u_riscv_cpu_inst_write_en),
    .stage2_flush(u_riscv_cpu_stage2_flush),
    .stage2_stall(u_riscv_cpu_stage2_stall),
    .stage1_valid_flush(u_riscv_cpu_stage1_valid_flush),
    .inst_ready_to_use(u_riscv_cpu_inst_ready_to_use),
    .inst_buffer_full(u_riscv_cpu_inst_buffer_full),
    .data_sram_en(u_riscv_cpu_data_sram_en),
    .data_sram_wen(u_riscv_cpu_data_sram_wen),
    .data_size(u_riscv_cpu_data_size),
    .data_sram_addr(u_riscv_cpu_data_sram_addr),
    .data_sram_wdata(u_riscv_cpu_data_sram_wdata),
    .data_cache(u_riscv_cpu_data_cache),
    .data_sram_rdata(u_riscv_cpu_data_sram_rdata),
    .data_stage2_stall(u_riscv_cpu_data_stage2_stall),
    .data_wstrb(u_riscv_cpu_data_wstrb),
    .data_fence_i_control(u_riscv_cpu_data_fence_i_control),
    .debug_wb_pc(u_riscv_cpu_debug_wb_pc),
    .debug_wb_rf_wen(u_riscv_cpu_debug_wb_rf_wen),
    .debug_wb_rf_wnum(u_riscv_cpu_debug_wb_rf_wnum),
    .debug_wb_rf_wdata(u_riscv_cpu_debug_wb_rf_wdata),
    .icache_tag_flush(u_riscv_cpu_icache_tag_flush)
  );
  inst_cache inst_cache ( // @[my_cpu_top.scala 128:30]
    .clock(inst_cache_clock),
    .reset(inst_cache_reset),
    .io_port_araddr(inst_cache_io_port_araddr),
    .io_port_arlen(inst_cache_io_port_arlen),
    .io_port_arburst(inst_cache_io_port_arburst),
    .io_port_arvalid(inst_cache_io_port_arvalid),
    .io_port_arready(inst_cache_io_port_arready),
    .io_port_rdata(inst_cache_io_port_rdata),
    .io_port_rlast(inst_cache_io_port_rlast),
    .io_port_rvalid(inst_cache_io_port_rvalid),
    .io_stage2_flush(inst_cache_io_stage2_flush),
    .io_stage2_stall(inst_cache_io_stage2_stall),
    .io_stage1_valid_flush(inst_cache_io_stage1_valid_flush),
    .io_inst_ready_to_use(inst_cache_io_inst_ready_to_use),
    .io_inst_buffer_full(inst_cache_io_inst_buffer_full),
    .io_v_addr_for_tlb(inst_cache_io_v_addr_for_tlb),
    .io_p_addr_for_tlb(inst_cache_io_p_addr_for_tlb),
    .io_sram_req(inst_cache_io_sram_req),
    .io_sram_addr(inst_cache_io_sram_addr),
    .io_sram_write_en(inst_cache_io_sram_write_en),
    .io_sram_rdata_L(inst_cache_io_sram_rdata_L),
    .io_sram_cache(inst_cache_io_sram_cache),
    .io_tag_valid_flush(inst_cache_io_tag_valid_flush)
  );
  data_cache data_cache ( // @[my_cpu_top.scala 130:30]
    .clock(data_cache_clock),
    .reset(data_cache_reset),
    .io_port_araddr(data_cache_io_port_araddr),
    .io_port_arlen(data_cache_io_port_arlen),
    .io_port_arsize(data_cache_io_port_arsize),
    .io_port_arburst(data_cache_io_port_arburst),
    .io_port_arvalid(data_cache_io_port_arvalid),
    .io_port_arready(data_cache_io_port_arready),
    .io_port_rdata(data_cache_io_port_rdata),
    .io_port_rlast(data_cache_io_port_rlast),
    .io_port_rvalid(data_cache_io_port_rvalid),
    .io_port_awaddr(data_cache_io_port_awaddr),
    .io_port_awlen(data_cache_io_port_awlen),
    .io_port_awsize(data_cache_io_port_awsize),
    .io_port_awburst(data_cache_io_port_awburst),
    .io_port_awvalid(data_cache_io_port_awvalid),
    .io_port_awready(data_cache_io_port_awready),
    .io_port_wdata(data_cache_io_port_wdata),
    .io_port_wstrb(data_cache_io_port_wstrb),
    .io_port_wlast(data_cache_io_port_wlast),
    .io_port_wvalid(data_cache_io_port_wvalid),
    .io_port_wready(data_cache_io_port_wready),
    .io_port_bvalid(data_cache_io_port_bvalid),
    .io_stage2_stall(data_cache_io_stage2_stall),
    .io_v_addr_for_tlb(data_cache_io_v_addr_for_tlb),
    .io_p_addr_for_tlb(data_cache_io_p_addr_for_tlb),
    .io_tlb_req(data_cache_io_tlb_req),
    .io_data_wstrb(data_cache_io_data_wstrb),
    .io_sram_req(data_cache_io_sram_req),
    .io_sram_wr(data_cache_io_sram_wr),
    .io_sram_size(data_cache_io_sram_size),
    .io_sram_addr(data_cache_io_sram_addr),
    .io_sram_wdata(data_cache_io_sram_wdata),
    .io_sram_rdata(data_cache_io_sram_rdata),
    .io_sram_cache(data_cache_io_sram_cache),
    .io_fence_i_control(data_cache_io_fence_i_control)
  );
  axi_cross_bar_addr_switch _axi_cross_bar ( // @[my_cpu_top.scala 132:32]
    .clock(_axi_cross_bar_clock),
    .reset(_axi_cross_bar_reset),
    .io_m_port_0_araddr(_axi_cross_bar_io_m_port_0_araddr),
    .io_m_port_0_arlen(_axi_cross_bar_io_m_port_0_arlen),
    .io_m_port_0_arburst(_axi_cross_bar_io_m_port_0_arburst),
    .io_m_port_0_arvalid(_axi_cross_bar_io_m_port_0_arvalid),
    .io_m_port_0_arready(_axi_cross_bar_io_m_port_0_arready),
    .io_m_port_0_rdata(_axi_cross_bar_io_m_port_0_rdata),
    .io_m_port_0_rlast(_axi_cross_bar_io_m_port_0_rlast),
    .io_m_port_0_rvalid(_axi_cross_bar_io_m_port_0_rvalid),
    .io_m_port_1_araddr(_axi_cross_bar_io_m_port_1_araddr),
    .io_m_port_1_arlen(_axi_cross_bar_io_m_port_1_arlen),
    .io_m_port_1_arsize(_axi_cross_bar_io_m_port_1_arsize),
    .io_m_port_1_arburst(_axi_cross_bar_io_m_port_1_arburst),
    .io_m_port_1_arvalid(_axi_cross_bar_io_m_port_1_arvalid),
    .io_m_port_1_arready(_axi_cross_bar_io_m_port_1_arready),
    .io_m_port_1_rdata(_axi_cross_bar_io_m_port_1_rdata),
    .io_m_port_1_rlast(_axi_cross_bar_io_m_port_1_rlast),
    .io_m_port_1_rvalid(_axi_cross_bar_io_m_port_1_rvalid),
    .io_m_port_1_awaddr(_axi_cross_bar_io_m_port_1_awaddr),
    .io_m_port_1_awlen(_axi_cross_bar_io_m_port_1_awlen),
    .io_m_port_1_awsize(_axi_cross_bar_io_m_port_1_awsize),
    .io_m_port_1_awburst(_axi_cross_bar_io_m_port_1_awburst),
    .io_m_port_1_awvalid(_axi_cross_bar_io_m_port_1_awvalid),
    .io_m_port_1_awready(_axi_cross_bar_io_m_port_1_awready),
    .io_m_port_1_wdata(_axi_cross_bar_io_m_port_1_wdata),
    .io_m_port_1_wstrb(_axi_cross_bar_io_m_port_1_wstrb),
    .io_m_port_1_wlast(_axi_cross_bar_io_m_port_1_wlast),
    .io_m_port_1_wvalid(_axi_cross_bar_io_m_port_1_wvalid),
    .io_m_port_1_wready(_axi_cross_bar_io_m_port_1_wready),
    .io_m_port_1_bvalid(_axi_cross_bar_io_m_port_1_bvalid),
    .io_s_port_0_arid(_axi_cross_bar_io_s_port_0_arid),
    .io_s_port_0_araddr(_axi_cross_bar_io_s_port_0_araddr),
    .io_s_port_0_arlen(_axi_cross_bar_io_s_port_0_arlen),
    .io_s_port_0_arsize(_axi_cross_bar_io_s_port_0_arsize),
    .io_s_port_0_arburst(_axi_cross_bar_io_s_port_0_arburst),
    .io_s_port_0_arvalid(_axi_cross_bar_io_s_port_0_arvalid),
    .io_s_port_0_arready(_axi_cross_bar_io_s_port_0_arready),
    .io_s_port_0_rdata(_axi_cross_bar_io_s_port_0_rdata),
    .io_s_port_0_rlast(_axi_cross_bar_io_s_port_0_rlast),
    .io_s_port_0_rvalid(_axi_cross_bar_io_s_port_0_rvalid),
    .io_s_port_0_rready(_axi_cross_bar_io_s_port_0_rready),
    .io_s_port_0_awid(_axi_cross_bar_io_s_port_0_awid),
    .io_s_port_0_awaddr(_axi_cross_bar_io_s_port_0_awaddr),
    .io_s_port_0_awlen(_axi_cross_bar_io_s_port_0_awlen),
    .io_s_port_0_awsize(_axi_cross_bar_io_s_port_0_awsize),
    .io_s_port_0_awburst(_axi_cross_bar_io_s_port_0_awburst),
    .io_s_port_0_awvalid(_axi_cross_bar_io_s_port_0_awvalid),
    .io_s_port_0_awready(_axi_cross_bar_io_s_port_0_awready),
    .io_s_port_0_wid(_axi_cross_bar_io_s_port_0_wid),
    .io_s_port_0_wdata(_axi_cross_bar_io_s_port_0_wdata),
    .io_s_port_0_wstrb(_axi_cross_bar_io_s_port_0_wstrb),
    .io_s_port_0_wlast(_axi_cross_bar_io_s_port_0_wlast),
    .io_s_port_0_wvalid(_axi_cross_bar_io_s_port_0_wvalid),
    .io_s_port_0_wready(_axi_cross_bar_io_s_port_0_wready),
    .io_s_port_0_bvalid(_axi_cross_bar_io_s_port_0_bvalid),
    .io_s_port_0_bready(_axi_cross_bar_io_s_port_0_bready),
    .io_s_port_1_araddr(_axi_cross_bar_io_s_port_1_araddr),
    .io_s_port_1_arvalid(_axi_cross_bar_io_s_port_1_arvalid),
    .io_s_port_1_rdata(_axi_cross_bar_io_s_port_1_rdata),
    .io_s_port_1_rlast(_axi_cross_bar_io_s_port_1_rlast),
    .io_s_port_1_rvalid(_axi_cross_bar_io_s_port_1_rvalid),
    .io_s_port_1_rready(_axi_cross_bar_io_s_port_1_rready),
    .io_s_port_1_awaddr(_axi_cross_bar_io_s_port_1_awaddr),
    .io_s_port_1_awsize(_axi_cross_bar_io_s_port_1_awsize),
    .io_s_port_1_awvalid(_axi_cross_bar_io_s_port_1_awvalid),
    .io_s_port_1_wdata(_axi_cross_bar_io_s_port_1_wdata),
    .io_s_port_1_wvalid(_axi_cross_bar_io_s_port_1_wvalid),
    .io_s_port_1_wready(_axi_cross_bar_io_s_port_1_wready),
    .io_s_port_1_bvalid(_axi_cross_bar_io_s_port_1_bvalid)
  );
  timer_periph timer_periph ( // @[my_cpu_top.scala 242:27]
    .clock(timer_periph_clock),
    .reset(timer_periph_reset),
    .io_axi_port_araddr(timer_periph_io_axi_port_araddr),
    .io_axi_port_arvalid(timer_periph_io_axi_port_arvalid),
    .io_axi_port_arready(timer_periph_io_axi_port_arready),
    .io_axi_port_rdata(timer_periph_io_axi_port_rdata),
    .io_axi_port_rlast(timer_periph_io_axi_port_rlast),
    .io_axi_port_rvalid(timer_periph_io_axi_port_rvalid),
    .io_axi_port_rready(timer_periph_io_axi_port_rready),
    .io_axi_port_awaddr(timer_periph_io_axi_port_awaddr),
    .io_axi_port_awsize(timer_periph_io_axi_port_awsize),
    .io_axi_port_awvalid(timer_periph_io_axi_port_awvalid),
    .io_axi_port_awready(timer_periph_io_axi_port_awready),
    .io_axi_port_wdata(timer_periph_io_axi_port_wdata),
    .io_axi_port_wvalid(timer_periph_io_axi_port_wvalid),
    .io_axi_port_wready(timer_periph_io_axi_port_wready),
    .io_axi_port_bvalid(timer_periph_io_axi_port_bvalid),
    .io_int_line(timer_periph_io_int_line)
  );
  assign axi_mem_port_arid = _axi_cross_bar_io_s_port_0_arid; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_araddr = _axi_cross_bar_io_s_port_0_araddr; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_arlen = _axi_cross_bar_io_s_port_0_arlen; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_arsize = _axi_cross_bar_io_s_port_0_arsize; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_arburst = _axi_cross_bar_io_s_port_0_arburst; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_arlock = 2'h0; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_arcache = 4'h0; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_arprot = 3'h0; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_arvalid = _axi_cross_bar_io_s_port_0_arvalid; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_rready = _axi_cross_bar_io_s_port_0_rready; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_awid = _axi_cross_bar_io_s_port_0_awid; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_awaddr = _axi_cross_bar_io_s_port_0_awaddr; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_awlen = _axi_cross_bar_io_s_port_0_awlen; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_awsize = _axi_cross_bar_io_s_port_0_awsize; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_awburst = _axi_cross_bar_io_s_port_0_awburst; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_awlock = 2'h0; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_awcache = 4'h0; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_awprot = 3'h0; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_awvalid = _axi_cross_bar_io_s_port_0_awvalid; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_wid = _axi_cross_bar_io_s_port_0_wid; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_wdata = _axi_cross_bar_io_s_port_0_wdata; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_wstrb = _axi_cross_bar_io_s_port_0_wstrb; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_wlast = _axi_cross_bar_io_s_port_0_wlast; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_wvalid = _axi_cross_bar_io_s_port_0_wvalid; // @[my_cpu_top.scala 236:18]
  assign axi_mem_port_bready = _axi_cross_bar_io_s_port_0_bready; // @[my_cpu_top.scala 236:18]
  assign debug_wb_pc = u_riscv_cpu_debug_wb_pc[31:0]; // @[my_cpu_top.scala 223:29]
  assign debug_wb_rf_wen = u_riscv_cpu_debug_wb_rf_wen; // @[my_cpu_top.scala 225:29]
  assign debug_wb_rf_wnum = u_riscv_cpu_debug_wb_rf_wnum; // @[my_cpu_top.scala 226:29]
  assign debug_wb_rf_wdata = u_riscv_cpu_debug_wb_rf_wdata[31:0]; // @[my_cpu_top.scala 224:29]
  assign u_riscv_cpu_ext_int_timer = timer_periph_io_int_line; // @[my_cpu_top.scala 245:31]
  assign u_riscv_cpu_resetn = aresetn; // @[my_cpu_top.scala 228:30]
  assign u_riscv_cpu_clk = aclk; // @[my_cpu_top.scala 227:30]
  assign u_riscv_cpu_inst_sram_rdata_L = inst_cache_io_sram_rdata_L; // @[my_cpu_top.scala 210:32]
  assign u_riscv_cpu_inst_write_en = inst_cache_io_sram_write_en; // @[my_cpu_top.scala 218:31]
  assign u_riscv_cpu_stage2_stall = inst_cache_io_stage2_stall; // @[my_cpu_top.scala 230:35]
  assign u_riscv_cpu_data_sram_rdata = data_cache_io_sram_rdata; // @[my_cpu_top.scala 197:28]
  assign u_riscv_cpu_data_stage2_stall = data_cache_io_stage2_stall; // @[my_cpu_top.scala 219:35]
  assign inst_cache_clock = aclk; // @[my_cpu_top.scala 124:23]
  assign inst_cache_reset = ~aresetn; // @[my_cpu_top.scala 124:42]
  assign inst_cache_io_port_arready = _axi_cross_bar_io_m_port_0_arready; // @[my_cpu_top.scala 238:33]
  assign inst_cache_io_port_rdata = _axi_cross_bar_io_m_port_0_rdata; // @[my_cpu_top.scala 238:33]
  assign inst_cache_io_port_rlast = _axi_cross_bar_io_m_port_0_rlast; // @[my_cpu_top.scala 238:33]
  assign inst_cache_io_port_rvalid = _axi_cross_bar_io_m_port_0_rvalid; // @[my_cpu_top.scala 238:33]
  assign inst_cache_io_stage2_flush = u_riscv_cpu_stage2_flush; // @[my_cpu_top.scala 233:31]
  assign inst_cache_io_stage1_valid_flush = u_riscv_cpu_stage1_valid_flush; // @[my_cpu_top.scala 351:37]
  assign inst_cache_io_inst_ready_to_use = u_riscv_cpu_inst_ready_to_use; // @[my_cpu_top.scala 352:36]
  assign inst_cache_io_inst_buffer_full = u_riscv_cpu_inst_buffer_full; // @[my_cpu_top.scala 353:37]
  assign inst_cache_io_p_addr_for_tlb = inst_cache_io_v_addr_for_tlb; // @[my_cpu_top.scala 168:38]
  assign inst_cache_io_sram_req = u_riscv_cpu_inst_sram_en; // @[my_cpu_top.scala 204:29]
  assign inst_cache_io_sram_addr = u_riscv_cpu_inst_sram_addr; // @[my_cpu_top.scala 201:29]
  assign inst_cache_io_sram_cache = u_riscv_cpu_inst_cache; // @[my_cpu_top.scala 203:29]
  assign inst_cache_io_tag_valid_flush = u_riscv_cpu_icache_tag_flush; // @[my_cpu_top.scala 234:34]
  assign data_cache_clock = aclk; // @[my_cpu_top.scala 124:23]
  assign data_cache_reset = ~aresetn; // @[my_cpu_top.scala 124:42]
  assign data_cache_io_port_arready = _axi_cross_bar_io_m_port_1_arready; // @[my_cpu_top.scala 239:33]
  assign data_cache_io_port_rdata = _axi_cross_bar_io_m_port_1_rdata; // @[my_cpu_top.scala 239:33]
  assign data_cache_io_port_rlast = _axi_cross_bar_io_m_port_1_rlast; // @[my_cpu_top.scala 239:33]
  assign data_cache_io_port_rvalid = _axi_cross_bar_io_m_port_1_rvalid; // @[my_cpu_top.scala 239:33]
  assign data_cache_io_port_awready = _axi_cross_bar_io_m_port_1_awready; // @[my_cpu_top.scala 239:33]
  assign data_cache_io_port_wready = _axi_cross_bar_io_m_port_1_wready; // @[my_cpu_top.scala 239:33]
  assign data_cache_io_port_bvalid = _axi_cross_bar_io_m_port_1_bvalid; // @[my_cpu_top.scala 239:33]
  assign data_cache_io_p_addr_for_tlb = data_cache_io_v_addr_for_tlb; // @[my_cpu_top.scala 169:38]
  assign data_cache_io_data_wstrb = u_riscv_cpu_data_wstrb; // @[my_cpu_top.scala 196:29]
  assign data_cache_io_sram_req = u_riscv_cpu_data_sram_en; // @[my_cpu_top.scala 192:23]
  assign data_cache_io_sram_wr = u_riscv_cpu_data_sram_wen; // @[my_cpu_top.scala 193:23]
  assign data_cache_io_sram_size = {{1'd0}, u_riscv_cpu_data_size}; // @[my_cpu_top.scala 190:22]
  assign data_cache_io_sram_addr = u_riscv_cpu_data_sram_addr; // @[my_cpu_top.scala 189:22]
  assign data_cache_io_sram_wdata = u_riscv_cpu_data_sram_wdata; // @[my_cpu_top.scala 194:23]
  assign data_cache_io_sram_cache = u_riscv_cpu_data_cache; // @[my_cpu_top.scala 191:23]
  assign data_cache_io_fence_i_control = u_riscv_cpu_data_fence_i_control; // @[my_cpu_top.scala 195:28]
  assign _axi_cross_bar_clock = aclk; // @[my_cpu_top.scala 124:23]
  assign _axi_cross_bar_reset = ~aresetn; // @[my_cpu_top.scala 124:42]
  assign _axi_cross_bar_io_m_port_0_araddr = inst_cache_io_port_araddr; // @[my_cpu_top.scala 238:33]
  assign _axi_cross_bar_io_m_port_0_arlen = inst_cache_io_port_arlen; // @[my_cpu_top.scala 238:33]
  assign _axi_cross_bar_io_m_port_0_arburst = inst_cache_io_port_arburst; // @[my_cpu_top.scala 238:33]
  assign _axi_cross_bar_io_m_port_0_arvalid = inst_cache_io_port_arvalid; // @[my_cpu_top.scala 238:33]
  assign _axi_cross_bar_io_m_port_1_araddr = data_cache_io_port_araddr; // @[my_cpu_top.scala 239:33]
  assign _axi_cross_bar_io_m_port_1_arlen = data_cache_io_port_arlen; // @[my_cpu_top.scala 239:33]
  assign _axi_cross_bar_io_m_port_1_arsize = data_cache_io_port_arsize; // @[my_cpu_top.scala 239:33]
  assign _axi_cross_bar_io_m_port_1_arburst = data_cache_io_port_arburst; // @[my_cpu_top.scala 239:33]
  assign _axi_cross_bar_io_m_port_1_arvalid = data_cache_io_port_arvalid; // @[my_cpu_top.scala 239:33]
  assign _axi_cross_bar_io_m_port_1_awaddr = data_cache_io_port_awaddr; // @[my_cpu_top.scala 239:33]
  assign _axi_cross_bar_io_m_port_1_awlen = data_cache_io_port_awlen; // @[my_cpu_top.scala 239:33]
  assign _axi_cross_bar_io_m_port_1_awsize = data_cache_io_port_awsize; // @[my_cpu_top.scala 239:33]
  assign _axi_cross_bar_io_m_port_1_awburst = data_cache_io_port_awburst; // @[my_cpu_top.scala 239:33]
  assign _axi_cross_bar_io_m_port_1_awvalid = data_cache_io_port_awvalid; // @[my_cpu_top.scala 239:33]
  assign _axi_cross_bar_io_m_port_1_wdata = data_cache_io_port_wdata; // @[my_cpu_top.scala 239:33]
  assign _axi_cross_bar_io_m_port_1_wstrb = data_cache_io_port_wstrb; // @[my_cpu_top.scala 239:33]
  assign _axi_cross_bar_io_m_port_1_wlast = data_cache_io_port_wlast; // @[my_cpu_top.scala 239:33]
  assign _axi_cross_bar_io_m_port_1_wvalid = data_cache_io_port_wvalid; // @[my_cpu_top.scala 239:33]
  assign _axi_cross_bar_io_s_port_0_arready = axi_mem_port_arready; // @[my_cpu_top.scala 236:18]
  assign _axi_cross_bar_io_s_port_0_rdata = axi_mem_port_rdata; // @[my_cpu_top.scala 236:18]
  assign _axi_cross_bar_io_s_port_0_rlast = axi_mem_port_rlast; // @[my_cpu_top.scala 236:18]
  assign _axi_cross_bar_io_s_port_0_rvalid = axi_mem_port_rvalid; // @[my_cpu_top.scala 236:18]
  assign _axi_cross_bar_io_s_port_0_awready = axi_mem_port_awready; // @[my_cpu_top.scala 236:18]
  assign _axi_cross_bar_io_s_port_0_wready = axi_mem_port_wready; // @[my_cpu_top.scala 236:18]
  assign _axi_cross_bar_io_s_port_0_bvalid = axi_mem_port_bvalid; // @[my_cpu_top.scala 236:18]
  assign _axi_cross_bar_io_s_port_1_rdata = timer_periph_io_axi_port_rdata; // @[my_cpu_top.scala 243:33]
  assign _axi_cross_bar_io_s_port_1_rlast = timer_periph_io_axi_port_rlast; // @[my_cpu_top.scala 243:33]
  assign _axi_cross_bar_io_s_port_1_rvalid = timer_periph_io_axi_port_rvalid; // @[my_cpu_top.scala 243:33]
  assign _axi_cross_bar_io_s_port_1_wready = timer_periph_io_axi_port_wready; // @[my_cpu_top.scala 243:33]
  assign _axi_cross_bar_io_s_port_1_bvalid = timer_periph_io_axi_port_bvalid; // @[my_cpu_top.scala 243:33]
  assign timer_periph_clock = aclk; // @[my_cpu_top.scala 124:23]
  assign timer_periph_reset = ~aresetn; // @[my_cpu_top.scala 124:42]
  assign timer_periph_io_axi_port_araddr = _axi_cross_bar_io_s_port_1_araddr; // @[my_cpu_top.scala 243:33]
  assign timer_periph_io_axi_port_arvalid = _axi_cross_bar_io_s_port_1_arvalid; // @[my_cpu_top.scala 243:33]
  assign timer_periph_io_axi_port_rready = _axi_cross_bar_io_s_port_1_rready; // @[my_cpu_top.scala 243:33]
  assign timer_periph_io_axi_port_awaddr = _axi_cross_bar_io_s_port_1_awaddr; // @[my_cpu_top.scala 243:33]
  assign timer_periph_io_axi_port_awsize = _axi_cross_bar_io_s_port_1_awsize; // @[my_cpu_top.scala 243:33]
  assign timer_periph_io_axi_port_awvalid = _axi_cross_bar_io_s_port_1_awvalid; // @[my_cpu_top.scala 243:33]
  assign timer_periph_io_axi_port_wdata = _axi_cross_bar_io_s_port_1_wdata; // @[my_cpu_top.scala 243:33]
  assign timer_periph_io_axi_port_wvalid = _axi_cross_bar_io_s_port_1_wvalid; // @[my_cpu_top.scala 243:33]
endmodule
