module Mux2(
  input   io_sel,
  input   io_in0,
  input   io_in1,
  output  io_out
);
  assign io_out = io_sel & io_in1 | ~io_sel & io_in0; // @[mux2.scala 15:33]
endmodule
module AND(
  input         clock,
  input         reset,
  input         io_a,
  input         io_d,
  input  [31:0] io_b,
  output        io_c,
  input         io_data_in,
  input  [6:0]  io_data_sel,
  output        io_data_out,
  output [31:0] io_out,
  input  [31:0] io_data_data_input,
  output [31:0] io_data_out_out_data_input
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
`endif // RANDOMIZE_REG_INIT
  wire  Mux2_test_io_sel; // @[AND.scala 30:25]
  wire  Mux2_test_io_in0; // @[AND.scala 30:25]
  wire  Mux2_test_io_in1; // @[AND.scala 30:25]
  wire  Mux2_test_io_out; // @[AND.scala 30:25]
  wire  Mux3_test_io_sel; // @[AND.scala 31:25]
  wire  Mux3_test_io_in0; // @[AND.scala 31:25]
  wire  Mux3_test_io_in1; // @[AND.scala 31:25]
  wire  Mux3_test_io_out; // @[AND.scala 31:25]
  wire  stage_decoder_pc_0_io_sel; // @[AND.scala 32:44]
  wire  stage_decoder_pc_0_io_in0; // @[AND.scala 32:44]
  wire  stage_decoder_pc_0_io_in1; // @[AND.scala 32:44]
  wire  stage_decoder_pc_0_io_out; // @[AND.scala 32:44]
  wire  stage_decoder_pc_1_io_sel; // @[AND.scala 32:44]
  wire  stage_decoder_pc_1_io_in0; // @[AND.scala 32:44]
  wire  stage_decoder_pc_1_io_in1; // @[AND.scala 32:44]
  wire  stage_decoder_pc_1_io_out; // @[AND.scala 32:44]
  reg [31:0] io_data_out_out_REG_data_input; // @[AND.scala 29:29]
  wire [1:0] _GEN_384 = {{1'd0}, io_a}; // @[Mux.scala 81:61]
  wire  _io_out_T_1 = stage_decoder_pc_0_io_out + stage_decoder_pc_1_io_out; // @[AND.scala 59:39]
  reg  lru_0; // @[AND.scala 61:20]
  reg  lru_1; // @[AND.scala 61:20]
  reg  lru_2; // @[AND.scala 61:20]
  reg  lru_3; // @[AND.scala 61:20]
  reg  lru_4; // @[AND.scala 61:20]
  reg  lru_5; // @[AND.scala 61:20]
  reg  lru_6; // @[AND.scala 61:20]
  reg  lru_7; // @[AND.scala 61:20]
  reg  lru_8; // @[AND.scala 61:20]
  reg  lru_9; // @[AND.scala 61:20]
  reg  lru_10; // @[AND.scala 61:20]
  reg  lru_11; // @[AND.scala 61:20]
  reg  lru_12; // @[AND.scala 61:20]
  reg  lru_13; // @[AND.scala 61:20]
  reg  lru_14; // @[AND.scala 61:20]
  reg  lru_15; // @[AND.scala 61:20]
  reg  lru_16; // @[AND.scala 61:20]
  reg  lru_17; // @[AND.scala 61:20]
  reg  lru_18; // @[AND.scala 61:20]
  reg  lru_19; // @[AND.scala 61:20]
  reg  lru_20; // @[AND.scala 61:20]
  reg  lru_21; // @[AND.scala 61:20]
  reg  lru_22; // @[AND.scala 61:20]
  reg  lru_23; // @[AND.scala 61:20]
  reg  lru_24; // @[AND.scala 61:20]
  reg  lru_25; // @[AND.scala 61:20]
  reg  lru_26; // @[AND.scala 61:20]
  reg  lru_27; // @[AND.scala 61:20]
  reg  lru_28; // @[AND.scala 61:20]
  reg  lru_29; // @[AND.scala 61:20]
  reg  lru_30; // @[AND.scala 61:20]
  reg  lru_31; // @[AND.scala 61:20]
  reg  lru_32; // @[AND.scala 61:20]
  reg  lru_33; // @[AND.scala 61:20]
  reg  lru_34; // @[AND.scala 61:20]
  reg  lru_35; // @[AND.scala 61:20]
  reg  lru_36; // @[AND.scala 61:20]
  reg  lru_37; // @[AND.scala 61:20]
  reg  lru_38; // @[AND.scala 61:20]
  reg  lru_39; // @[AND.scala 61:20]
  reg  lru_40; // @[AND.scala 61:20]
  reg  lru_41; // @[AND.scala 61:20]
  reg  lru_42; // @[AND.scala 61:20]
  reg  lru_43; // @[AND.scala 61:20]
  reg  lru_44; // @[AND.scala 61:20]
  reg  lru_45; // @[AND.scala 61:20]
  reg  lru_46; // @[AND.scala 61:20]
  reg  lru_47; // @[AND.scala 61:20]
  reg  lru_48; // @[AND.scala 61:20]
  reg  lru_49; // @[AND.scala 61:20]
  reg  lru_50; // @[AND.scala 61:20]
  reg  lru_51; // @[AND.scala 61:20]
  reg  lru_52; // @[AND.scala 61:20]
  reg  lru_53; // @[AND.scala 61:20]
  reg  lru_54; // @[AND.scala 61:20]
  reg  lru_55; // @[AND.scala 61:20]
  reg  lru_56; // @[AND.scala 61:20]
  reg  lru_57; // @[AND.scala 61:20]
  reg  lru_58; // @[AND.scala 61:20]
  reg  lru_59; // @[AND.scala 61:20]
  reg  lru_60; // @[AND.scala 61:20]
  reg  lru_61; // @[AND.scala 61:20]
  reg  lru_62; // @[AND.scala 61:20]
  reg  lru_63; // @[AND.scala 61:20]
  reg  lru_64; // @[AND.scala 61:20]
  reg  lru_65; // @[AND.scala 61:20]
  reg  lru_66; // @[AND.scala 61:20]
  reg  lru_67; // @[AND.scala 61:20]
  reg  lru_68; // @[AND.scala 61:20]
  reg  lru_69; // @[AND.scala 61:20]
  reg  lru_70; // @[AND.scala 61:20]
  reg  lru_71; // @[AND.scala 61:20]
  reg  lru_72; // @[AND.scala 61:20]
  reg  lru_73; // @[AND.scala 61:20]
  reg  lru_74; // @[AND.scala 61:20]
  reg  lru_75; // @[AND.scala 61:20]
  reg  lru_76; // @[AND.scala 61:20]
  reg  lru_77; // @[AND.scala 61:20]
  reg  lru_78; // @[AND.scala 61:20]
  reg  lru_79; // @[AND.scala 61:20]
  reg  lru_80; // @[AND.scala 61:20]
  reg  lru_81; // @[AND.scala 61:20]
  reg  lru_82; // @[AND.scala 61:20]
  reg  lru_83; // @[AND.scala 61:20]
  reg  lru_84; // @[AND.scala 61:20]
  reg  lru_85; // @[AND.scala 61:20]
  reg  lru_86; // @[AND.scala 61:20]
  reg  lru_87; // @[AND.scala 61:20]
  reg  lru_88; // @[AND.scala 61:20]
  reg  lru_89; // @[AND.scala 61:20]
  reg  lru_90; // @[AND.scala 61:20]
  reg  lru_91; // @[AND.scala 61:20]
  reg  lru_92; // @[AND.scala 61:20]
  reg  lru_93; // @[AND.scala 61:20]
  reg  lru_94; // @[AND.scala 61:20]
  reg  lru_95; // @[AND.scala 61:20]
  reg  lru_96; // @[AND.scala 61:20]
  reg  lru_97; // @[AND.scala 61:20]
  reg  lru_98; // @[AND.scala 61:20]
  reg  lru_99; // @[AND.scala 61:20]
  reg  lru_100; // @[AND.scala 61:20]
  reg  lru_101; // @[AND.scala 61:20]
  reg  lru_102; // @[AND.scala 61:20]
  reg  lru_103; // @[AND.scala 61:20]
  reg  lru_104; // @[AND.scala 61:20]
  reg  lru_105; // @[AND.scala 61:20]
  reg  lru_106; // @[AND.scala 61:20]
  reg  lru_107; // @[AND.scala 61:20]
  reg  lru_108; // @[AND.scala 61:20]
  reg  lru_109; // @[AND.scala 61:20]
  reg  lru_110; // @[AND.scala 61:20]
  reg  lru_111; // @[AND.scala 61:20]
  reg  lru_112; // @[AND.scala 61:20]
  reg  lru_113; // @[AND.scala 61:20]
  reg  lru_114; // @[AND.scala 61:20]
  reg  lru_115; // @[AND.scala 61:20]
  reg  lru_116; // @[AND.scala 61:20]
  reg  lru_117; // @[AND.scala 61:20]
  reg  lru_118; // @[AND.scala 61:20]
  reg  lru_119; // @[AND.scala 61:20]
  reg  lru_120; // @[AND.scala 61:20]
  reg  lru_121; // @[AND.scala 61:20]
  reg  lru_122; // @[AND.scala 61:20]
  reg  lru_123; // @[AND.scala 61:20]
  reg  lru_124; // @[AND.scala 61:20]
  reg  lru_125; // @[AND.scala 61:20]
  reg  lru_126; // @[AND.scala 61:20]
  reg  lru_127; // @[AND.scala 61:20]
  wire [6:0] _io_data_out_T_2 = {1'h0,io_data_sel[5:0]}; // @[Cat.scala 31:58]
  wire [7:0] _io_data_out_T_3 = {1'h1,io_data_sel}; // @[Cat.scala 31:58]
  wire  _GEN_129 = 7'h1 == _io_data_out_T_2 ? lru_1 : lru_0; // @[AND.scala 63:{21,21}]
  wire  _GEN_130 = 7'h2 == _io_data_out_T_2 ? lru_2 : _GEN_129; // @[AND.scala 63:{21,21}]
  wire  _GEN_131 = 7'h3 == _io_data_out_T_2 ? lru_3 : _GEN_130; // @[AND.scala 63:{21,21}]
  wire  _GEN_132 = 7'h4 == _io_data_out_T_2 ? lru_4 : _GEN_131; // @[AND.scala 63:{21,21}]
  wire  _GEN_133 = 7'h5 == _io_data_out_T_2 ? lru_5 : _GEN_132; // @[AND.scala 63:{21,21}]
  wire  _GEN_134 = 7'h6 == _io_data_out_T_2 ? lru_6 : _GEN_133; // @[AND.scala 63:{21,21}]
  wire  _GEN_135 = 7'h7 == _io_data_out_T_2 ? lru_7 : _GEN_134; // @[AND.scala 63:{21,21}]
  wire  _GEN_136 = 7'h8 == _io_data_out_T_2 ? lru_8 : _GEN_135; // @[AND.scala 63:{21,21}]
  wire  _GEN_137 = 7'h9 == _io_data_out_T_2 ? lru_9 : _GEN_136; // @[AND.scala 63:{21,21}]
  wire  _GEN_138 = 7'ha == _io_data_out_T_2 ? lru_10 : _GEN_137; // @[AND.scala 63:{21,21}]
  wire  _GEN_139 = 7'hb == _io_data_out_T_2 ? lru_11 : _GEN_138; // @[AND.scala 63:{21,21}]
  wire  _GEN_140 = 7'hc == _io_data_out_T_2 ? lru_12 : _GEN_139; // @[AND.scala 63:{21,21}]
  wire  _GEN_141 = 7'hd == _io_data_out_T_2 ? lru_13 : _GEN_140; // @[AND.scala 63:{21,21}]
  wire  _GEN_142 = 7'he == _io_data_out_T_2 ? lru_14 : _GEN_141; // @[AND.scala 63:{21,21}]
  wire  _GEN_143 = 7'hf == _io_data_out_T_2 ? lru_15 : _GEN_142; // @[AND.scala 63:{21,21}]
  wire  _GEN_144 = 7'h10 == _io_data_out_T_2 ? lru_16 : _GEN_143; // @[AND.scala 63:{21,21}]
  wire  _GEN_145 = 7'h11 == _io_data_out_T_2 ? lru_17 : _GEN_144; // @[AND.scala 63:{21,21}]
  wire  _GEN_146 = 7'h12 == _io_data_out_T_2 ? lru_18 : _GEN_145; // @[AND.scala 63:{21,21}]
  wire  _GEN_147 = 7'h13 == _io_data_out_T_2 ? lru_19 : _GEN_146; // @[AND.scala 63:{21,21}]
  wire  _GEN_148 = 7'h14 == _io_data_out_T_2 ? lru_20 : _GEN_147; // @[AND.scala 63:{21,21}]
  wire  _GEN_149 = 7'h15 == _io_data_out_T_2 ? lru_21 : _GEN_148; // @[AND.scala 63:{21,21}]
  wire  _GEN_150 = 7'h16 == _io_data_out_T_2 ? lru_22 : _GEN_149; // @[AND.scala 63:{21,21}]
  wire  _GEN_151 = 7'h17 == _io_data_out_T_2 ? lru_23 : _GEN_150; // @[AND.scala 63:{21,21}]
  wire  _GEN_152 = 7'h18 == _io_data_out_T_2 ? lru_24 : _GEN_151; // @[AND.scala 63:{21,21}]
  wire  _GEN_153 = 7'h19 == _io_data_out_T_2 ? lru_25 : _GEN_152; // @[AND.scala 63:{21,21}]
  wire  _GEN_154 = 7'h1a == _io_data_out_T_2 ? lru_26 : _GEN_153; // @[AND.scala 63:{21,21}]
  wire  _GEN_155 = 7'h1b == _io_data_out_T_2 ? lru_27 : _GEN_154; // @[AND.scala 63:{21,21}]
  wire  _GEN_156 = 7'h1c == _io_data_out_T_2 ? lru_28 : _GEN_155; // @[AND.scala 63:{21,21}]
  wire  _GEN_157 = 7'h1d == _io_data_out_T_2 ? lru_29 : _GEN_156; // @[AND.scala 63:{21,21}]
  wire  _GEN_158 = 7'h1e == _io_data_out_T_2 ? lru_30 : _GEN_157; // @[AND.scala 63:{21,21}]
  wire  _GEN_159 = 7'h1f == _io_data_out_T_2 ? lru_31 : _GEN_158; // @[AND.scala 63:{21,21}]
  wire  _GEN_160 = 7'h20 == _io_data_out_T_2 ? lru_32 : _GEN_159; // @[AND.scala 63:{21,21}]
  wire  _GEN_161 = 7'h21 == _io_data_out_T_2 ? lru_33 : _GEN_160; // @[AND.scala 63:{21,21}]
  wire  _GEN_162 = 7'h22 == _io_data_out_T_2 ? lru_34 : _GEN_161; // @[AND.scala 63:{21,21}]
  wire  _GEN_163 = 7'h23 == _io_data_out_T_2 ? lru_35 : _GEN_162; // @[AND.scala 63:{21,21}]
  wire  _GEN_164 = 7'h24 == _io_data_out_T_2 ? lru_36 : _GEN_163; // @[AND.scala 63:{21,21}]
  wire  _GEN_165 = 7'h25 == _io_data_out_T_2 ? lru_37 : _GEN_164; // @[AND.scala 63:{21,21}]
  wire  _GEN_166 = 7'h26 == _io_data_out_T_2 ? lru_38 : _GEN_165; // @[AND.scala 63:{21,21}]
  wire  _GEN_167 = 7'h27 == _io_data_out_T_2 ? lru_39 : _GEN_166; // @[AND.scala 63:{21,21}]
  wire  _GEN_168 = 7'h28 == _io_data_out_T_2 ? lru_40 : _GEN_167; // @[AND.scala 63:{21,21}]
  wire  _GEN_169 = 7'h29 == _io_data_out_T_2 ? lru_41 : _GEN_168; // @[AND.scala 63:{21,21}]
  wire  _GEN_170 = 7'h2a == _io_data_out_T_2 ? lru_42 : _GEN_169; // @[AND.scala 63:{21,21}]
  wire  _GEN_171 = 7'h2b == _io_data_out_T_2 ? lru_43 : _GEN_170; // @[AND.scala 63:{21,21}]
  wire  _GEN_172 = 7'h2c == _io_data_out_T_2 ? lru_44 : _GEN_171; // @[AND.scala 63:{21,21}]
  wire  _GEN_173 = 7'h2d == _io_data_out_T_2 ? lru_45 : _GEN_172; // @[AND.scala 63:{21,21}]
  wire  _GEN_174 = 7'h2e == _io_data_out_T_2 ? lru_46 : _GEN_173; // @[AND.scala 63:{21,21}]
  wire  _GEN_175 = 7'h2f == _io_data_out_T_2 ? lru_47 : _GEN_174; // @[AND.scala 63:{21,21}]
  wire  _GEN_176 = 7'h30 == _io_data_out_T_2 ? lru_48 : _GEN_175; // @[AND.scala 63:{21,21}]
  wire  _GEN_177 = 7'h31 == _io_data_out_T_2 ? lru_49 : _GEN_176; // @[AND.scala 63:{21,21}]
  wire  _GEN_178 = 7'h32 == _io_data_out_T_2 ? lru_50 : _GEN_177; // @[AND.scala 63:{21,21}]
  wire  _GEN_179 = 7'h33 == _io_data_out_T_2 ? lru_51 : _GEN_178; // @[AND.scala 63:{21,21}]
  wire  _GEN_180 = 7'h34 == _io_data_out_T_2 ? lru_52 : _GEN_179; // @[AND.scala 63:{21,21}]
  wire  _GEN_181 = 7'h35 == _io_data_out_T_2 ? lru_53 : _GEN_180; // @[AND.scala 63:{21,21}]
  wire  _GEN_182 = 7'h36 == _io_data_out_T_2 ? lru_54 : _GEN_181; // @[AND.scala 63:{21,21}]
  wire  _GEN_183 = 7'h37 == _io_data_out_T_2 ? lru_55 : _GEN_182; // @[AND.scala 63:{21,21}]
  wire  _GEN_184 = 7'h38 == _io_data_out_T_2 ? lru_56 : _GEN_183; // @[AND.scala 63:{21,21}]
  wire  _GEN_185 = 7'h39 == _io_data_out_T_2 ? lru_57 : _GEN_184; // @[AND.scala 63:{21,21}]
  wire  _GEN_186 = 7'h3a == _io_data_out_T_2 ? lru_58 : _GEN_185; // @[AND.scala 63:{21,21}]
  wire  _GEN_187 = 7'h3b == _io_data_out_T_2 ? lru_59 : _GEN_186; // @[AND.scala 63:{21,21}]
  wire  _GEN_188 = 7'h3c == _io_data_out_T_2 ? lru_60 : _GEN_187; // @[AND.scala 63:{21,21}]
  wire  _GEN_189 = 7'h3d == _io_data_out_T_2 ? lru_61 : _GEN_188; // @[AND.scala 63:{21,21}]
  wire  _GEN_190 = 7'h3e == _io_data_out_T_2 ? lru_62 : _GEN_189; // @[AND.scala 63:{21,21}]
  wire  _GEN_191 = 7'h3f == _io_data_out_T_2 ? lru_63 : _GEN_190; // @[AND.scala 63:{21,21}]
  wire  _GEN_192 = 7'h40 == _io_data_out_T_2 ? lru_64 : _GEN_191; // @[AND.scala 63:{21,21}]
  wire  _GEN_193 = 7'h41 == _io_data_out_T_2 ? lru_65 : _GEN_192; // @[AND.scala 63:{21,21}]
  wire  _GEN_194 = 7'h42 == _io_data_out_T_2 ? lru_66 : _GEN_193; // @[AND.scala 63:{21,21}]
  wire  _GEN_195 = 7'h43 == _io_data_out_T_2 ? lru_67 : _GEN_194; // @[AND.scala 63:{21,21}]
  wire  _GEN_196 = 7'h44 == _io_data_out_T_2 ? lru_68 : _GEN_195; // @[AND.scala 63:{21,21}]
  wire  _GEN_197 = 7'h45 == _io_data_out_T_2 ? lru_69 : _GEN_196; // @[AND.scala 63:{21,21}]
  wire  _GEN_198 = 7'h46 == _io_data_out_T_2 ? lru_70 : _GEN_197; // @[AND.scala 63:{21,21}]
  wire  _GEN_199 = 7'h47 == _io_data_out_T_2 ? lru_71 : _GEN_198; // @[AND.scala 63:{21,21}]
  wire  _GEN_200 = 7'h48 == _io_data_out_T_2 ? lru_72 : _GEN_199; // @[AND.scala 63:{21,21}]
  wire  _GEN_201 = 7'h49 == _io_data_out_T_2 ? lru_73 : _GEN_200; // @[AND.scala 63:{21,21}]
  wire  _GEN_202 = 7'h4a == _io_data_out_T_2 ? lru_74 : _GEN_201; // @[AND.scala 63:{21,21}]
  wire  _GEN_203 = 7'h4b == _io_data_out_T_2 ? lru_75 : _GEN_202; // @[AND.scala 63:{21,21}]
  wire  _GEN_204 = 7'h4c == _io_data_out_T_2 ? lru_76 : _GEN_203; // @[AND.scala 63:{21,21}]
  wire  _GEN_205 = 7'h4d == _io_data_out_T_2 ? lru_77 : _GEN_204; // @[AND.scala 63:{21,21}]
  wire  _GEN_206 = 7'h4e == _io_data_out_T_2 ? lru_78 : _GEN_205; // @[AND.scala 63:{21,21}]
  wire  _GEN_207 = 7'h4f == _io_data_out_T_2 ? lru_79 : _GEN_206; // @[AND.scala 63:{21,21}]
  wire  _GEN_208 = 7'h50 == _io_data_out_T_2 ? lru_80 : _GEN_207; // @[AND.scala 63:{21,21}]
  wire  _GEN_209 = 7'h51 == _io_data_out_T_2 ? lru_81 : _GEN_208; // @[AND.scala 63:{21,21}]
  wire  _GEN_210 = 7'h52 == _io_data_out_T_2 ? lru_82 : _GEN_209; // @[AND.scala 63:{21,21}]
  wire  _GEN_211 = 7'h53 == _io_data_out_T_2 ? lru_83 : _GEN_210; // @[AND.scala 63:{21,21}]
  wire  _GEN_212 = 7'h54 == _io_data_out_T_2 ? lru_84 : _GEN_211; // @[AND.scala 63:{21,21}]
  wire  _GEN_213 = 7'h55 == _io_data_out_T_2 ? lru_85 : _GEN_212; // @[AND.scala 63:{21,21}]
  wire  _GEN_214 = 7'h56 == _io_data_out_T_2 ? lru_86 : _GEN_213; // @[AND.scala 63:{21,21}]
  wire  _GEN_215 = 7'h57 == _io_data_out_T_2 ? lru_87 : _GEN_214; // @[AND.scala 63:{21,21}]
  wire  _GEN_216 = 7'h58 == _io_data_out_T_2 ? lru_88 : _GEN_215; // @[AND.scala 63:{21,21}]
  wire  _GEN_217 = 7'h59 == _io_data_out_T_2 ? lru_89 : _GEN_216; // @[AND.scala 63:{21,21}]
  wire  _GEN_218 = 7'h5a == _io_data_out_T_2 ? lru_90 : _GEN_217; // @[AND.scala 63:{21,21}]
  wire  _GEN_219 = 7'h5b == _io_data_out_T_2 ? lru_91 : _GEN_218; // @[AND.scala 63:{21,21}]
  wire  _GEN_220 = 7'h5c == _io_data_out_T_2 ? lru_92 : _GEN_219; // @[AND.scala 63:{21,21}]
  wire  _GEN_221 = 7'h5d == _io_data_out_T_2 ? lru_93 : _GEN_220; // @[AND.scala 63:{21,21}]
  wire  _GEN_222 = 7'h5e == _io_data_out_T_2 ? lru_94 : _GEN_221; // @[AND.scala 63:{21,21}]
  wire  _GEN_223 = 7'h5f == _io_data_out_T_2 ? lru_95 : _GEN_222; // @[AND.scala 63:{21,21}]
  wire  _GEN_224 = 7'h60 == _io_data_out_T_2 ? lru_96 : _GEN_223; // @[AND.scala 63:{21,21}]
  wire  _GEN_225 = 7'h61 == _io_data_out_T_2 ? lru_97 : _GEN_224; // @[AND.scala 63:{21,21}]
  wire  _GEN_226 = 7'h62 == _io_data_out_T_2 ? lru_98 : _GEN_225; // @[AND.scala 63:{21,21}]
  wire  _GEN_227 = 7'h63 == _io_data_out_T_2 ? lru_99 : _GEN_226; // @[AND.scala 63:{21,21}]
  wire  _GEN_228 = 7'h64 == _io_data_out_T_2 ? lru_100 : _GEN_227; // @[AND.scala 63:{21,21}]
  wire  _GEN_229 = 7'h65 == _io_data_out_T_2 ? lru_101 : _GEN_228; // @[AND.scala 63:{21,21}]
  wire  _GEN_230 = 7'h66 == _io_data_out_T_2 ? lru_102 : _GEN_229; // @[AND.scala 63:{21,21}]
  wire  _GEN_231 = 7'h67 == _io_data_out_T_2 ? lru_103 : _GEN_230; // @[AND.scala 63:{21,21}]
  wire  _GEN_232 = 7'h68 == _io_data_out_T_2 ? lru_104 : _GEN_231; // @[AND.scala 63:{21,21}]
  wire  _GEN_233 = 7'h69 == _io_data_out_T_2 ? lru_105 : _GEN_232; // @[AND.scala 63:{21,21}]
  wire  _GEN_234 = 7'h6a == _io_data_out_T_2 ? lru_106 : _GEN_233; // @[AND.scala 63:{21,21}]
  wire  _GEN_235 = 7'h6b == _io_data_out_T_2 ? lru_107 : _GEN_234; // @[AND.scala 63:{21,21}]
  wire  _GEN_236 = 7'h6c == _io_data_out_T_2 ? lru_108 : _GEN_235; // @[AND.scala 63:{21,21}]
  wire  _GEN_237 = 7'h6d == _io_data_out_T_2 ? lru_109 : _GEN_236; // @[AND.scala 63:{21,21}]
  wire  _GEN_238 = 7'h6e == _io_data_out_T_2 ? lru_110 : _GEN_237; // @[AND.scala 63:{21,21}]
  wire  _GEN_239 = 7'h6f == _io_data_out_T_2 ? lru_111 : _GEN_238; // @[AND.scala 63:{21,21}]
  wire  _GEN_240 = 7'h70 == _io_data_out_T_2 ? lru_112 : _GEN_239; // @[AND.scala 63:{21,21}]
  wire  _GEN_241 = 7'h71 == _io_data_out_T_2 ? lru_113 : _GEN_240; // @[AND.scala 63:{21,21}]
  wire  _GEN_242 = 7'h72 == _io_data_out_T_2 ? lru_114 : _GEN_241; // @[AND.scala 63:{21,21}]
  wire  _GEN_243 = 7'h73 == _io_data_out_T_2 ? lru_115 : _GEN_242; // @[AND.scala 63:{21,21}]
  wire  _GEN_244 = 7'h74 == _io_data_out_T_2 ? lru_116 : _GEN_243; // @[AND.scala 63:{21,21}]
  wire  _GEN_245 = 7'h75 == _io_data_out_T_2 ? lru_117 : _GEN_244; // @[AND.scala 63:{21,21}]
  wire  _GEN_246 = 7'h76 == _io_data_out_T_2 ? lru_118 : _GEN_245; // @[AND.scala 63:{21,21}]
  wire  _GEN_247 = 7'h77 == _io_data_out_T_2 ? lru_119 : _GEN_246; // @[AND.scala 63:{21,21}]
  wire  _GEN_248 = 7'h78 == _io_data_out_T_2 ? lru_120 : _GEN_247; // @[AND.scala 63:{21,21}]
  wire  _GEN_249 = 7'h79 == _io_data_out_T_2 ? lru_121 : _GEN_248; // @[AND.scala 63:{21,21}]
  wire  _GEN_250 = 7'h7a == _io_data_out_T_2 ? lru_122 : _GEN_249; // @[AND.scala 63:{21,21}]
  wire  _GEN_251 = 7'h7b == _io_data_out_T_2 ? lru_123 : _GEN_250; // @[AND.scala 63:{21,21}]
  wire  _GEN_252 = 7'h7c == _io_data_out_T_2 ? lru_124 : _GEN_251; // @[AND.scala 63:{21,21}]
  wire  _GEN_253 = 7'h7d == _io_data_out_T_2 ? lru_125 : _GEN_252; // @[AND.scala 63:{21,21}]
  wire  _GEN_254 = 7'h7e == _io_data_out_T_2 ? lru_126 : _GEN_253; // @[AND.scala 63:{21,21}]
  wire  _GEN_255 = 7'h7f == _io_data_out_T_2 ? lru_127 : _GEN_254; // @[AND.scala 63:{21,21}]
  wire  _GEN_257 = 7'h1 == _io_data_out_T_3[6:0] ? lru_1 : lru_0; // @[AND.scala 63:{21,21}]
  wire  _GEN_258 = 7'h2 == _io_data_out_T_3[6:0] ? lru_2 : _GEN_257; // @[AND.scala 63:{21,21}]
  wire  _GEN_259 = 7'h3 == _io_data_out_T_3[6:0] ? lru_3 : _GEN_258; // @[AND.scala 63:{21,21}]
  wire  _GEN_260 = 7'h4 == _io_data_out_T_3[6:0] ? lru_4 : _GEN_259; // @[AND.scala 63:{21,21}]
  wire  _GEN_261 = 7'h5 == _io_data_out_T_3[6:0] ? lru_5 : _GEN_260; // @[AND.scala 63:{21,21}]
  wire  _GEN_262 = 7'h6 == _io_data_out_T_3[6:0] ? lru_6 : _GEN_261; // @[AND.scala 63:{21,21}]
  wire  _GEN_263 = 7'h7 == _io_data_out_T_3[6:0] ? lru_7 : _GEN_262; // @[AND.scala 63:{21,21}]
  wire  _GEN_264 = 7'h8 == _io_data_out_T_3[6:0] ? lru_8 : _GEN_263; // @[AND.scala 63:{21,21}]
  wire  _GEN_265 = 7'h9 == _io_data_out_T_3[6:0] ? lru_9 : _GEN_264; // @[AND.scala 63:{21,21}]
  wire  _GEN_266 = 7'ha == _io_data_out_T_3[6:0] ? lru_10 : _GEN_265; // @[AND.scala 63:{21,21}]
  wire  _GEN_267 = 7'hb == _io_data_out_T_3[6:0] ? lru_11 : _GEN_266; // @[AND.scala 63:{21,21}]
  wire  _GEN_268 = 7'hc == _io_data_out_T_3[6:0] ? lru_12 : _GEN_267; // @[AND.scala 63:{21,21}]
  wire  _GEN_269 = 7'hd == _io_data_out_T_3[6:0] ? lru_13 : _GEN_268; // @[AND.scala 63:{21,21}]
  wire  _GEN_270 = 7'he == _io_data_out_T_3[6:0] ? lru_14 : _GEN_269; // @[AND.scala 63:{21,21}]
  wire  _GEN_271 = 7'hf == _io_data_out_T_3[6:0] ? lru_15 : _GEN_270; // @[AND.scala 63:{21,21}]
  wire  _GEN_272 = 7'h10 == _io_data_out_T_3[6:0] ? lru_16 : _GEN_271; // @[AND.scala 63:{21,21}]
  wire  _GEN_273 = 7'h11 == _io_data_out_T_3[6:0] ? lru_17 : _GEN_272; // @[AND.scala 63:{21,21}]
  wire  _GEN_274 = 7'h12 == _io_data_out_T_3[6:0] ? lru_18 : _GEN_273; // @[AND.scala 63:{21,21}]
  wire  _GEN_275 = 7'h13 == _io_data_out_T_3[6:0] ? lru_19 : _GEN_274; // @[AND.scala 63:{21,21}]
  wire  _GEN_276 = 7'h14 == _io_data_out_T_3[6:0] ? lru_20 : _GEN_275; // @[AND.scala 63:{21,21}]
  wire  _GEN_277 = 7'h15 == _io_data_out_T_3[6:0] ? lru_21 : _GEN_276; // @[AND.scala 63:{21,21}]
  wire  _GEN_278 = 7'h16 == _io_data_out_T_3[6:0] ? lru_22 : _GEN_277; // @[AND.scala 63:{21,21}]
  wire  _GEN_279 = 7'h17 == _io_data_out_T_3[6:0] ? lru_23 : _GEN_278; // @[AND.scala 63:{21,21}]
  wire  _GEN_280 = 7'h18 == _io_data_out_T_3[6:0] ? lru_24 : _GEN_279; // @[AND.scala 63:{21,21}]
  wire  _GEN_281 = 7'h19 == _io_data_out_T_3[6:0] ? lru_25 : _GEN_280; // @[AND.scala 63:{21,21}]
  wire  _GEN_282 = 7'h1a == _io_data_out_T_3[6:0] ? lru_26 : _GEN_281; // @[AND.scala 63:{21,21}]
  wire  _GEN_283 = 7'h1b == _io_data_out_T_3[6:0] ? lru_27 : _GEN_282; // @[AND.scala 63:{21,21}]
  wire  _GEN_284 = 7'h1c == _io_data_out_T_3[6:0] ? lru_28 : _GEN_283; // @[AND.scala 63:{21,21}]
  wire  _GEN_285 = 7'h1d == _io_data_out_T_3[6:0] ? lru_29 : _GEN_284; // @[AND.scala 63:{21,21}]
  wire  _GEN_286 = 7'h1e == _io_data_out_T_3[6:0] ? lru_30 : _GEN_285; // @[AND.scala 63:{21,21}]
  wire  _GEN_287 = 7'h1f == _io_data_out_T_3[6:0] ? lru_31 : _GEN_286; // @[AND.scala 63:{21,21}]
  wire  _GEN_288 = 7'h20 == _io_data_out_T_3[6:0] ? lru_32 : _GEN_287; // @[AND.scala 63:{21,21}]
  wire  _GEN_289 = 7'h21 == _io_data_out_T_3[6:0] ? lru_33 : _GEN_288; // @[AND.scala 63:{21,21}]
  wire  _GEN_290 = 7'h22 == _io_data_out_T_3[6:0] ? lru_34 : _GEN_289; // @[AND.scala 63:{21,21}]
  wire  _GEN_291 = 7'h23 == _io_data_out_T_3[6:0] ? lru_35 : _GEN_290; // @[AND.scala 63:{21,21}]
  wire  _GEN_292 = 7'h24 == _io_data_out_T_3[6:0] ? lru_36 : _GEN_291; // @[AND.scala 63:{21,21}]
  wire  _GEN_293 = 7'h25 == _io_data_out_T_3[6:0] ? lru_37 : _GEN_292; // @[AND.scala 63:{21,21}]
  wire  _GEN_294 = 7'h26 == _io_data_out_T_3[6:0] ? lru_38 : _GEN_293; // @[AND.scala 63:{21,21}]
  wire  _GEN_295 = 7'h27 == _io_data_out_T_3[6:0] ? lru_39 : _GEN_294; // @[AND.scala 63:{21,21}]
  wire  _GEN_296 = 7'h28 == _io_data_out_T_3[6:0] ? lru_40 : _GEN_295; // @[AND.scala 63:{21,21}]
  wire  _GEN_297 = 7'h29 == _io_data_out_T_3[6:0] ? lru_41 : _GEN_296; // @[AND.scala 63:{21,21}]
  wire  _GEN_298 = 7'h2a == _io_data_out_T_3[6:0] ? lru_42 : _GEN_297; // @[AND.scala 63:{21,21}]
  wire  _GEN_299 = 7'h2b == _io_data_out_T_3[6:0] ? lru_43 : _GEN_298; // @[AND.scala 63:{21,21}]
  wire  _GEN_300 = 7'h2c == _io_data_out_T_3[6:0] ? lru_44 : _GEN_299; // @[AND.scala 63:{21,21}]
  wire  _GEN_301 = 7'h2d == _io_data_out_T_3[6:0] ? lru_45 : _GEN_300; // @[AND.scala 63:{21,21}]
  wire  _GEN_302 = 7'h2e == _io_data_out_T_3[6:0] ? lru_46 : _GEN_301; // @[AND.scala 63:{21,21}]
  wire  _GEN_303 = 7'h2f == _io_data_out_T_3[6:0] ? lru_47 : _GEN_302; // @[AND.scala 63:{21,21}]
  wire  _GEN_304 = 7'h30 == _io_data_out_T_3[6:0] ? lru_48 : _GEN_303; // @[AND.scala 63:{21,21}]
  wire  _GEN_305 = 7'h31 == _io_data_out_T_3[6:0] ? lru_49 : _GEN_304; // @[AND.scala 63:{21,21}]
  wire  _GEN_306 = 7'h32 == _io_data_out_T_3[6:0] ? lru_50 : _GEN_305; // @[AND.scala 63:{21,21}]
  wire  _GEN_307 = 7'h33 == _io_data_out_T_3[6:0] ? lru_51 : _GEN_306; // @[AND.scala 63:{21,21}]
  wire  _GEN_308 = 7'h34 == _io_data_out_T_3[6:0] ? lru_52 : _GEN_307; // @[AND.scala 63:{21,21}]
  wire  _GEN_309 = 7'h35 == _io_data_out_T_3[6:0] ? lru_53 : _GEN_308; // @[AND.scala 63:{21,21}]
  wire  _GEN_310 = 7'h36 == _io_data_out_T_3[6:0] ? lru_54 : _GEN_309; // @[AND.scala 63:{21,21}]
  wire  _GEN_311 = 7'h37 == _io_data_out_T_3[6:0] ? lru_55 : _GEN_310; // @[AND.scala 63:{21,21}]
  wire  _GEN_312 = 7'h38 == _io_data_out_T_3[6:0] ? lru_56 : _GEN_311; // @[AND.scala 63:{21,21}]
  wire  _GEN_313 = 7'h39 == _io_data_out_T_3[6:0] ? lru_57 : _GEN_312; // @[AND.scala 63:{21,21}]
  wire  _GEN_314 = 7'h3a == _io_data_out_T_3[6:0] ? lru_58 : _GEN_313; // @[AND.scala 63:{21,21}]
  wire  _GEN_315 = 7'h3b == _io_data_out_T_3[6:0] ? lru_59 : _GEN_314; // @[AND.scala 63:{21,21}]
  wire  _GEN_316 = 7'h3c == _io_data_out_T_3[6:0] ? lru_60 : _GEN_315; // @[AND.scala 63:{21,21}]
  wire  _GEN_317 = 7'h3d == _io_data_out_T_3[6:0] ? lru_61 : _GEN_316; // @[AND.scala 63:{21,21}]
  wire  _GEN_318 = 7'h3e == _io_data_out_T_3[6:0] ? lru_62 : _GEN_317; // @[AND.scala 63:{21,21}]
  wire  _GEN_319 = 7'h3f == _io_data_out_T_3[6:0] ? lru_63 : _GEN_318; // @[AND.scala 63:{21,21}]
  wire  _GEN_320 = 7'h40 == _io_data_out_T_3[6:0] ? lru_64 : _GEN_319; // @[AND.scala 63:{21,21}]
  wire  _GEN_321 = 7'h41 == _io_data_out_T_3[6:0] ? lru_65 : _GEN_320; // @[AND.scala 63:{21,21}]
  wire  _GEN_322 = 7'h42 == _io_data_out_T_3[6:0] ? lru_66 : _GEN_321; // @[AND.scala 63:{21,21}]
  wire  _GEN_323 = 7'h43 == _io_data_out_T_3[6:0] ? lru_67 : _GEN_322; // @[AND.scala 63:{21,21}]
  wire  _GEN_324 = 7'h44 == _io_data_out_T_3[6:0] ? lru_68 : _GEN_323; // @[AND.scala 63:{21,21}]
  wire  _GEN_325 = 7'h45 == _io_data_out_T_3[6:0] ? lru_69 : _GEN_324; // @[AND.scala 63:{21,21}]
  wire  _GEN_326 = 7'h46 == _io_data_out_T_3[6:0] ? lru_70 : _GEN_325; // @[AND.scala 63:{21,21}]
  wire  _GEN_327 = 7'h47 == _io_data_out_T_3[6:0] ? lru_71 : _GEN_326; // @[AND.scala 63:{21,21}]
  wire  _GEN_328 = 7'h48 == _io_data_out_T_3[6:0] ? lru_72 : _GEN_327; // @[AND.scala 63:{21,21}]
  wire  _GEN_329 = 7'h49 == _io_data_out_T_3[6:0] ? lru_73 : _GEN_328; // @[AND.scala 63:{21,21}]
  wire  _GEN_330 = 7'h4a == _io_data_out_T_3[6:0] ? lru_74 : _GEN_329; // @[AND.scala 63:{21,21}]
  wire  _GEN_331 = 7'h4b == _io_data_out_T_3[6:0] ? lru_75 : _GEN_330; // @[AND.scala 63:{21,21}]
  wire  _GEN_332 = 7'h4c == _io_data_out_T_3[6:0] ? lru_76 : _GEN_331; // @[AND.scala 63:{21,21}]
  wire  _GEN_333 = 7'h4d == _io_data_out_T_3[6:0] ? lru_77 : _GEN_332; // @[AND.scala 63:{21,21}]
  wire  _GEN_334 = 7'h4e == _io_data_out_T_3[6:0] ? lru_78 : _GEN_333; // @[AND.scala 63:{21,21}]
  wire  _GEN_335 = 7'h4f == _io_data_out_T_3[6:0] ? lru_79 : _GEN_334; // @[AND.scala 63:{21,21}]
  wire  _GEN_336 = 7'h50 == _io_data_out_T_3[6:0] ? lru_80 : _GEN_335; // @[AND.scala 63:{21,21}]
  wire  _GEN_337 = 7'h51 == _io_data_out_T_3[6:0] ? lru_81 : _GEN_336; // @[AND.scala 63:{21,21}]
  wire  _GEN_338 = 7'h52 == _io_data_out_T_3[6:0] ? lru_82 : _GEN_337; // @[AND.scala 63:{21,21}]
  wire  _GEN_339 = 7'h53 == _io_data_out_T_3[6:0] ? lru_83 : _GEN_338; // @[AND.scala 63:{21,21}]
  wire  _GEN_340 = 7'h54 == _io_data_out_T_3[6:0] ? lru_84 : _GEN_339; // @[AND.scala 63:{21,21}]
  wire  _GEN_341 = 7'h55 == _io_data_out_T_3[6:0] ? lru_85 : _GEN_340; // @[AND.scala 63:{21,21}]
  wire  _GEN_342 = 7'h56 == _io_data_out_T_3[6:0] ? lru_86 : _GEN_341; // @[AND.scala 63:{21,21}]
  wire  _GEN_343 = 7'h57 == _io_data_out_T_3[6:0] ? lru_87 : _GEN_342; // @[AND.scala 63:{21,21}]
  wire  _GEN_344 = 7'h58 == _io_data_out_T_3[6:0] ? lru_88 : _GEN_343; // @[AND.scala 63:{21,21}]
  wire  _GEN_345 = 7'h59 == _io_data_out_T_3[6:0] ? lru_89 : _GEN_344; // @[AND.scala 63:{21,21}]
  wire  _GEN_346 = 7'h5a == _io_data_out_T_3[6:0] ? lru_90 : _GEN_345; // @[AND.scala 63:{21,21}]
  wire  _GEN_347 = 7'h5b == _io_data_out_T_3[6:0] ? lru_91 : _GEN_346; // @[AND.scala 63:{21,21}]
  wire  _GEN_348 = 7'h5c == _io_data_out_T_3[6:0] ? lru_92 : _GEN_347; // @[AND.scala 63:{21,21}]
  wire  _GEN_349 = 7'h5d == _io_data_out_T_3[6:0] ? lru_93 : _GEN_348; // @[AND.scala 63:{21,21}]
  wire  _GEN_350 = 7'h5e == _io_data_out_T_3[6:0] ? lru_94 : _GEN_349; // @[AND.scala 63:{21,21}]
  wire  _GEN_351 = 7'h5f == _io_data_out_T_3[6:0] ? lru_95 : _GEN_350; // @[AND.scala 63:{21,21}]
  wire  _GEN_352 = 7'h60 == _io_data_out_T_3[6:0] ? lru_96 : _GEN_351; // @[AND.scala 63:{21,21}]
  wire  _GEN_353 = 7'h61 == _io_data_out_T_3[6:0] ? lru_97 : _GEN_352; // @[AND.scala 63:{21,21}]
  wire  _GEN_354 = 7'h62 == _io_data_out_T_3[6:0] ? lru_98 : _GEN_353; // @[AND.scala 63:{21,21}]
  wire  _GEN_355 = 7'h63 == _io_data_out_T_3[6:0] ? lru_99 : _GEN_354; // @[AND.scala 63:{21,21}]
  wire  _GEN_356 = 7'h64 == _io_data_out_T_3[6:0] ? lru_100 : _GEN_355; // @[AND.scala 63:{21,21}]
  wire  _GEN_357 = 7'h65 == _io_data_out_T_3[6:0] ? lru_101 : _GEN_356; // @[AND.scala 63:{21,21}]
  wire  _GEN_358 = 7'h66 == _io_data_out_T_3[6:0] ? lru_102 : _GEN_357; // @[AND.scala 63:{21,21}]
  wire  _GEN_359 = 7'h67 == _io_data_out_T_3[6:0] ? lru_103 : _GEN_358; // @[AND.scala 63:{21,21}]
  wire  _GEN_360 = 7'h68 == _io_data_out_T_3[6:0] ? lru_104 : _GEN_359; // @[AND.scala 63:{21,21}]
  wire  _GEN_361 = 7'h69 == _io_data_out_T_3[6:0] ? lru_105 : _GEN_360; // @[AND.scala 63:{21,21}]
  wire  _GEN_362 = 7'h6a == _io_data_out_T_3[6:0] ? lru_106 : _GEN_361; // @[AND.scala 63:{21,21}]
  wire  _GEN_363 = 7'h6b == _io_data_out_T_3[6:0] ? lru_107 : _GEN_362; // @[AND.scala 63:{21,21}]
  wire  _GEN_364 = 7'h6c == _io_data_out_T_3[6:0] ? lru_108 : _GEN_363; // @[AND.scala 63:{21,21}]
  wire  _GEN_365 = 7'h6d == _io_data_out_T_3[6:0] ? lru_109 : _GEN_364; // @[AND.scala 63:{21,21}]
  wire  _GEN_366 = 7'h6e == _io_data_out_T_3[6:0] ? lru_110 : _GEN_365; // @[AND.scala 63:{21,21}]
  wire  _GEN_367 = 7'h6f == _io_data_out_T_3[6:0] ? lru_111 : _GEN_366; // @[AND.scala 63:{21,21}]
  wire  _GEN_368 = 7'h70 == _io_data_out_T_3[6:0] ? lru_112 : _GEN_367; // @[AND.scala 63:{21,21}]
  wire  _GEN_369 = 7'h71 == _io_data_out_T_3[6:0] ? lru_113 : _GEN_368; // @[AND.scala 63:{21,21}]
  wire  _GEN_370 = 7'h72 == _io_data_out_T_3[6:0] ? lru_114 : _GEN_369; // @[AND.scala 63:{21,21}]
  wire  _GEN_371 = 7'h73 == _io_data_out_T_3[6:0] ? lru_115 : _GEN_370; // @[AND.scala 63:{21,21}]
  wire  _GEN_372 = 7'h74 == _io_data_out_T_3[6:0] ? lru_116 : _GEN_371; // @[AND.scala 63:{21,21}]
  wire  _GEN_373 = 7'h75 == _io_data_out_T_3[6:0] ? lru_117 : _GEN_372; // @[AND.scala 63:{21,21}]
  wire  _GEN_374 = 7'h76 == _io_data_out_T_3[6:0] ? lru_118 : _GEN_373; // @[AND.scala 63:{21,21}]
  wire  _GEN_375 = 7'h77 == _io_data_out_T_3[6:0] ? lru_119 : _GEN_374; // @[AND.scala 63:{21,21}]
  wire  _GEN_376 = 7'h78 == _io_data_out_T_3[6:0] ? lru_120 : _GEN_375; // @[AND.scala 63:{21,21}]
  wire  _GEN_377 = 7'h79 == _io_data_out_T_3[6:0] ? lru_121 : _GEN_376; // @[AND.scala 63:{21,21}]
  wire  _GEN_378 = 7'h7a == _io_data_out_T_3[6:0] ? lru_122 : _GEN_377; // @[AND.scala 63:{21,21}]
  wire  _GEN_379 = 7'h7b == _io_data_out_T_3[6:0] ? lru_123 : _GEN_378; // @[AND.scala 63:{21,21}]
  wire  _GEN_380 = 7'h7c == _io_data_out_T_3[6:0] ? lru_124 : _GEN_379; // @[AND.scala 63:{21,21}]
  wire  _GEN_381 = 7'h7d == _io_data_out_T_3[6:0] ? lru_125 : _GEN_380; // @[AND.scala 63:{21,21}]
  wire  _GEN_382 = 7'h7e == _io_data_out_T_3[6:0] ? lru_126 : _GEN_381; // @[AND.scala 63:{21,21}]
  wire  _GEN_383 = 7'h7f == _io_data_out_T_3[6:0] ? lru_127 : _GEN_382; // @[AND.scala 63:{21,21}]
  Mux2 Mux2_test ( // @[AND.scala 30:25]
    .io_sel(Mux2_test_io_sel),
    .io_in0(Mux2_test_io_in0),
    .io_in1(Mux2_test_io_in1),
    .io_out(Mux2_test_io_out)
  );
  Mux2 Mux3_test ( // @[AND.scala 31:25]
    .io_sel(Mux3_test_io_sel),
    .io_in0(Mux3_test_io_in0),
    .io_in1(Mux3_test_io_in1),
    .io_out(Mux3_test_io_out)
  );
  Mux2 stage_decoder_pc_0 ( // @[AND.scala 32:44]
    .io_sel(stage_decoder_pc_0_io_sel),
    .io_in0(stage_decoder_pc_0_io_in0),
    .io_in1(stage_decoder_pc_0_io_in1),
    .io_out(stage_decoder_pc_0_io_out)
  );
  Mux2 stage_decoder_pc_1 ( // @[AND.scala 32:44]
    .io_sel(stage_decoder_pc_1_io_sel),
    .io_in0(stage_decoder_pc_1_io_in0),
    .io_in1(stage_decoder_pc_1_io_in1),
    .io_out(stage_decoder_pc_1_io_out)
  );
  assign io_c = 2'h3 == _GEN_384 ? stage_decoder_pc_1_io_out : io_a & stage_decoder_pc_0_io_out; // @[Mux.scala 81:58]
  assign io_data_out = io_data_sel[6] ? _GEN_255 : _GEN_383; // @[AND.scala 63:21]
  assign io_out = {{31'd0}, _io_out_T_1}; // @[AND.scala 59:10]
  assign io_data_out_out_data_input = io_data_out_out_REG_data_input; // @[AND.scala 29:19]
  assign Mux2_test_io_sel = io_d; // @[AND.scala 43:20]
  assign Mux2_test_io_in0 = io_a; // @[AND.scala 41:20]
  assign Mux2_test_io_in1 = io_b[0]; // @[AND.scala 42:20]
  assign Mux3_test_io_sel = Mux2_test_io_sel; // @[AND.scala 47:20]
  assign Mux3_test_io_in0 = Mux2_test_io_in0; // @[AND.scala 45:20]
  assign Mux3_test_io_in1 = Mux2_test_io_in1; // @[AND.scala 46:20]
  assign stage_decoder_pc_0_io_sel = io_d; // @[AND.scala 52:32]
  assign stage_decoder_pc_0_io_in0 = io_a; // @[AND.scala 50:32]
  assign stage_decoder_pc_0_io_in1 = io_b[0]; // @[AND.scala 51:32]
  assign stage_decoder_pc_1_io_sel = io_d; // @[AND.scala 52:32]
  assign stage_decoder_pc_1_io_in0 = io_a; // @[AND.scala 50:32]
  assign stage_decoder_pc_1_io_in1 = io_b[0]; // @[AND.scala 51:32]
  always @(posedge clock) begin
    io_data_out_out_REG_data_input <= io_data_data_input; // @[AND.scala 29:29]
    if (reset) begin // @[AND.scala 61:20]
      lru_0 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h0 == io_data_sel) begin // @[AND.scala 62:20]
      lru_0 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_1 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h1 == io_data_sel) begin // @[AND.scala 62:20]
      lru_1 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_2 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h2 == io_data_sel) begin // @[AND.scala 62:20]
      lru_2 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_3 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h3 == io_data_sel) begin // @[AND.scala 62:20]
      lru_3 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_4 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h4 == io_data_sel) begin // @[AND.scala 62:20]
      lru_4 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_5 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h5 == io_data_sel) begin // @[AND.scala 62:20]
      lru_5 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_6 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h6 == io_data_sel) begin // @[AND.scala 62:20]
      lru_6 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_7 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h7 == io_data_sel) begin // @[AND.scala 62:20]
      lru_7 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_8 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h8 == io_data_sel) begin // @[AND.scala 62:20]
      lru_8 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_9 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h9 == io_data_sel) begin // @[AND.scala 62:20]
      lru_9 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_10 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'ha == io_data_sel) begin // @[AND.scala 62:20]
      lru_10 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_11 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'hb == io_data_sel) begin // @[AND.scala 62:20]
      lru_11 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_12 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'hc == io_data_sel) begin // @[AND.scala 62:20]
      lru_12 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_13 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'hd == io_data_sel) begin // @[AND.scala 62:20]
      lru_13 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_14 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'he == io_data_sel) begin // @[AND.scala 62:20]
      lru_14 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_15 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'hf == io_data_sel) begin // @[AND.scala 62:20]
      lru_15 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_16 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h10 == io_data_sel) begin // @[AND.scala 62:20]
      lru_16 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_17 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h11 == io_data_sel) begin // @[AND.scala 62:20]
      lru_17 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_18 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h12 == io_data_sel) begin // @[AND.scala 62:20]
      lru_18 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_19 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h13 == io_data_sel) begin // @[AND.scala 62:20]
      lru_19 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_20 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h14 == io_data_sel) begin // @[AND.scala 62:20]
      lru_20 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_21 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h15 == io_data_sel) begin // @[AND.scala 62:20]
      lru_21 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_22 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h16 == io_data_sel) begin // @[AND.scala 62:20]
      lru_22 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_23 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h17 == io_data_sel) begin // @[AND.scala 62:20]
      lru_23 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_24 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h18 == io_data_sel) begin // @[AND.scala 62:20]
      lru_24 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_25 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h19 == io_data_sel) begin // @[AND.scala 62:20]
      lru_25 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_26 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h1a == io_data_sel) begin // @[AND.scala 62:20]
      lru_26 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_27 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h1b == io_data_sel) begin // @[AND.scala 62:20]
      lru_27 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_28 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h1c == io_data_sel) begin // @[AND.scala 62:20]
      lru_28 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_29 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h1d == io_data_sel) begin // @[AND.scala 62:20]
      lru_29 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_30 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h1e == io_data_sel) begin // @[AND.scala 62:20]
      lru_30 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_31 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h1f == io_data_sel) begin // @[AND.scala 62:20]
      lru_31 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_32 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h20 == io_data_sel) begin // @[AND.scala 62:20]
      lru_32 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_33 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h21 == io_data_sel) begin // @[AND.scala 62:20]
      lru_33 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_34 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h22 == io_data_sel) begin // @[AND.scala 62:20]
      lru_34 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_35 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h23 == io_data_sel) begin // @[AND.scala 62:20]
      lru_35 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_36 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h24 == io_data_sel) begin // @[AND.scala 62:20]
      lru_36 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_37 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h25 == io_data_sel) begin // @[AND.scala 62:20]
      lru_37 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_38 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h26 == io_data_sel) begin // @[AND.scala 62:20]
      lru_38 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_39 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h27 == io_data_sel) begin // @[AND.scala 62:20]
      lru_39 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_40 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h28 == io_data_sel) begin // @[AND.scala 62:20]
      lru_40 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_41 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h29 == io_data_sel) begin // @[AND.scala 62:20]
      lru_41 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_42 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h2a == io_data_sel) begin // @[AND.scala 62:20]
      lru_42 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_43 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h2b == io_data_sel) begin // @[AND.scala 62:20]
      lru_43 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_44 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h2c == io_data_sel) begin // @[AND.scala 62:20]
      lru_44 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_45 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h2d == io_data_sel) begin // @[AND.scala 62:20]
      lru_45 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_46 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h2e == io_data_sel) begin // @[AND.scala 62:20]
      lru_46 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_47 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h2f == io_data_sel) begin // @[AND.scala 62:20]
      lru_47 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_48 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h30 == io_data_sel) begin // @[AND.scala 62:20]
      lru_48 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_49 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h31 == io_data_sel) begin // @[AND.scala 62:20]
      lru_49 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_50 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h32 == io_data_sel) begin // @[AND.scala 62:20]
      lru_50 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_51 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h33 == io_data_sel) begin // @[AND.scala 62:20]
      lru_51 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_52 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h34 == io_data_sel) begin // @[AND.scala 62:20]
      lru_52 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_53 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h35 == io_data_sel) begin // @[AND.scala 62:20]
      lru_53 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_54 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h36 == io_data_sel) begin // @[AND.scala 62:20]
      lru_54 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_55 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h37 == io_data_sel) begin // @[AND.scala 62:20]
      lru_55 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_56 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h38 == io_data_sel) begin // @[AND.scala 62:20]
      lru_56 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_57 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h39 == io_data_sel) begin // @[AND.scala 62:20]
      lru_57 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_58 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h3a == io_data_sel) begin // @[AND.scala 62:20]
      lru_58 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_59 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h3b == io_data_sel) begin // @[AND.scala 62:20]
      lru_59 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_60 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h3c == io_data_sel) begin // @[AND.scala 62:20]
      lru_60 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_61 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h3d == io_data_sel) begin // @[AND.scala 62:20]
      lru_61 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_62 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h3e == io_data_sel) begin // @[AND.scala 62:20]
      lru_62 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_63 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h3f == io_data_sel) begin // @[AND.scala 62:20]
      lru_63 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_64 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h40 == io_data_sel) begin // @[AND.scala 62:20]
      lru_64 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_65 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h41 == io_data_sel) begin // @[AND.scala 62:20]
      lru_65 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_66 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h42 == io_data_sel) begin // @[AND.scala 62:20]
      lru_66 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_67 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h43 == io_data_sel) begin // @[AND.scala 62:20]
      lru_67 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_68 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h44 == io_data_sel) begin // @[AND.scala 62:20]
      lru_68 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_69 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h45 == io_data_sel) begin // @[AND.scala 62:20]
      lru_69 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_70 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h46 == io_data_sel) begin // @[AND.scala 62:20]
      lru_70 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_71 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h47 == io_data_sel) begin // @[AND.scala 62:20]
      lru_71 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_72 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h48 == io_data_sel) begin // @[AND.scala 62:20]
      lru_72 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_73 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h49 == io_data_sel) begin // @[AND.scala 62:20]
      lru_73 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_74 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h4a == io_data_sel) begin // @[AND.scala 62:20]
      lru_74 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_75 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h4b == io_data_sel) begin // @[AND.scala 62:20]
      lru_75 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_76 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h4c == io_data_sel) begin // @[AND.scala 62:20]
      lru_76 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_77 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h4d == io_data_sel) begin // @[AND.scala 62:20]
      lru_77 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_78 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h4e == io_data_sel) begin // @[AND.scala 62:20]
      lru_78 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_79 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h4f == io_data_sel) begin // @[AND.scala 62:20]
      lru_79 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_80 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h50 == io_data_sel) begin // @[AND.scala 62:20]
      lru_80 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_81 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h51 == io_data_sel) begin // @[AND.scala 62:20]
      lru_81 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_82 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h52 == io_data_sel) begin // @[AND.scala 62:20]
      lru_82 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_83 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h53 == io_data_sel) begin // @[AND.scala 62:20]
      lru_83 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_84 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h54 == io_data_sel) begin // @[AND.scala 62:20]
      lru_84 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_85 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h55 == io_data_sel) begin // @[AND.scala 62:20]
      lru_85 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_86 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h56 == io_data_sel) begin // @[AND.scala 62:20]
      lru_86 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_87 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h57 == io_data_sel) begin // @[AND.scala 62:20]
      lru_87 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_88 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h58 == io_data_sel) begin // @[AND.scala 62:20]
      lru_88 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_89 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h59 == io_data_sel) begin // @[AND.scala 62:20]
      lru_89 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_90 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h5a == io_data_sel) begin // @[AND.scala 62:20]
      lru_90 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_91 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h5b == io_data_sel) begin // @[AND.scala 62:20]
      lru_91 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_92 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h5c == io_data_sel) begin // @[AND.scala 62:20]
      lru_92 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_93 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h5d == io_data_sel) begin // @[AND.scala 62:20]
      lru_93 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_94 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h5e == io_data_sel) begin // @[AND.scala 62:20]
      lru_94 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_95 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h5f == io_data_sel) begin // @[AND.scala 62:20]
      lru_95 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_96 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h60 == io_data_sel) begin // @[AND.scala 62:20]
      lru_96 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_97 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h61 == io_data_sel) begin // @[AND.scala 62:20]
      lru_97 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_98 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h62 == io_data_sel) begin // @[AND.scala 62:20]
      lru_98 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_99 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h63 == io_data_sel) begin // @[AND.scala 62:20]
      lru_99 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_100 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h64 == io_data_sel) begin // @[AND.scala 62:20]
      lru_100 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_101 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h65 == io_data_sel) begin // @[AND.scala 62:20]
      lru_101 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_102 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h66 == io_data_sel) begin // @[AND.scala 62:20]
      lru_102 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_103 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h67 == io_data_sel) begin // @[AND.scala 62:20]
      lru_103 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_104 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h68 == io_data_sel) begin // @[AND.scala 62:20]
      lru_104 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_105 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h69 == io_data_sel) begin // @[AND.scala 62:20]
      lru_105 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_106 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h6a == io_data_sel) begin // @[AND.scala 62:20]
      lru_106 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_107 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h6b == io_data_sel) begin // @[AND.scala 62:20]
      lru_107 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_108 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h6c == io_data_sel) begin // @[AND.scala 62:20]
      lru_108 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_109 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h6d == io_data_sel) begin // @[AND.scala 62:20]
      lru_109 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_110 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h6e == io_data_sel) begin // @[AND.scala 62:20]
      lru_110 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_111 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h6f == io_data_sel) begin // @[AND.scala 62:20]
      lru_111 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_112 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h70 == io_data_sel) begin // @[AND.scala 62:20]
      lru_112 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_113 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h71 == io_data_sel) begin // @[AND.scala 62:20]
      lru_113 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_114 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h72 == io_data_sel) begin // @[AND.scala 62:20]
      lru_114 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_115 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h73 == io_data_sel) begin // @[AND.scala 62:20]
      lru_115 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_116 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h74 == io_data_sel) begin // @[AND.scala 62:20]
      lru_116 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_117 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h75 == io_data_sel) begin // @[AND.scala 62:20]
      lru_117 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_118 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h76 == io_data_sel) begin // @[AND.scala 62:20]
      lru_118 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_119 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h77 == io_data_sel) begin // @[AND.scala 62:20]
      lru_119 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_120 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h78 == io_data_sel) begin // @[AND.scala 62:20]
      lru_120 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_121 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h79 == io_data_sel) begin // @[AND.scala 62:20]
      lru_121 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_122 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h7a == io_data_sel) begin // @[AND.scala 62:20]
      lru_122 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_123 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h7b == io_data_sel) begin // @[AND.scala 62:20]
      lru_123 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_124 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h7c == io_data_sel) begin // @[AND.scala 62:20]
      lru_124 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_125 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h7d == io_data_sel) begin // @[AND.scala 62:20]
      lru_125 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_126 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h7e == io_data_sel) begin // @[AND.scala 62:20]
      lru_126 <= io_data_in; // @[AND.scala 62:20]
    end
    if (reset) begin // @[AND.scala 61:20]
      lru_127 <= 1'h0; // @[AND.scala 61:20]
    end else if (7'h7f == io_data_sel) begin // @[AND.scala 62:20]
      lru_127 <= io_data_in; // @[AND.scala 62:20]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_data_out_out_REG_data_input = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  lru_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  lru_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  lru_2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  lru_3 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  lru_4 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  lru_5 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  lru_6 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  lru_7 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  lru_8 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  lru_9 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  lru_10 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  lru_11 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  lru_12 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  lru_13 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  lru_14 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  lru_15 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  lru_16 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  lru_17 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  lru_18 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  lru_19 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  lru_20 = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  lru_21 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  lru_22 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  lru_23 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  lru_24 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  lru_25 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  lru_26 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  lru_27 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  lru_28 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  lru_29 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  lru_30 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  lru_31 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  lru_32 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  lru_33 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  lru_34 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  lru_35 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  lru_36 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  lru_37 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  lru_38 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  lru_39 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  lru_40 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  lru_41 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  lru_42 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  lru_43 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  lru_44 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  lru_45 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  lru_46 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  lru_47 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  lru_48 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  lru_49 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  lru_50 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  lru_51 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  lru_52 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  lru_53 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  lru_54 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  lru_55 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  lru_56 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  lru_57 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  lru_58 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  lru_59 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  lru_60 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  lru_61 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  lru_62 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  lru_63 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  lru_64 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  lru_65 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  lru_66 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  lru_67 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  lru_68 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  lru_69 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  lru_70 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  lru_71 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  lru_72 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  lru_73 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  lru_74 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  lru_75 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  lru_76 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  lru_77 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  lru_78 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  lru_79 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  lru_80 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  lru_81 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  lru_82 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  lru_83 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  lru_84 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  lru_85 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  lru_86 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  lru_87 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  lru_88 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  lru_89 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  lru_90 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  lru_91 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  lru_92 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  lru_93 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  lru_94 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  lru_95 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  lru_96 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  lru_97 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  lru_98 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  lru_99 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  lru_100 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  lru_101 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  lru_102 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  lru_103 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  lru_104 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  lru_105 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  lru_106 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  lru_107 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  lru_108 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  lru_109 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  lru_110 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  lru_111 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  lru_112 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  lru_113 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  lru_114 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  lru_115 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  lru_116 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  lru_117 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  lru_118 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  lru_119 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  lru_120 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  lru_121 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  lru_122 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  lru_123 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  lru_124 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  lru_125 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  lru_126 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  lru_127 = _RAND_128[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
